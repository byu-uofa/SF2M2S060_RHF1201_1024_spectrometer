
--+----------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.numeric_STD.all;

entity DataCtrl is
  --+----------
  -- Generic declarations
  --+----------
  generic(
          DataVecSize_g   :integer := 56;
          WdVecSize_g     :integer := 16;
          ByteSize_g      :integer := 8;
          NibbleSize_g    :integer := 4
      );

  --+----------
  -- Port name declarations
  --+----------
  port   (
       CLK100     :in  std_logic;
       RST        :in  std_logic;
       
       ADC_CLK_1  :out std_logic;
       ADC_CLK_2  :out std_logic; 
       
       ADC_D1_d   :in  std_logic_vector(11 downto 0); /* synthesis preserve=1*/
       ADC_DR1_d  :in  std_logic; /* synthesis preserve=1*/
               
       ADC_D2_d   :in  std_logic_vector(11 downto 0); /* synthesis preserve=1*/   
       ADC_DR2_d  :in  std_logic; /* synthesis preserve=1*/
       
       PEAK_FL_C1 :out  std_logic;

       
       i_PEAK_THD          :in std_logic_vector(11 downto 0);
       i_PEAK_THD_pos      :in std_logic_vector(11 downto 0);
       
       i_DR1_EN            : in std_logic;
       i_DR2_EN            : in std_logic;
       
       PEAK_C1             :out std_logic_vector(WdVecSize_g-5 downto 0);
       PEAK_C2             :out std_logic_vector(WdVecSize_g-5 downto 0);
       
       
       TIMESTAMP_C1          :out  std_logic_vector(DataVecSize_g-WdVecSize_g-1 downto 0);
       TIMESTAMP_C2          :out  std_logic_vector(DataVecSize_g-WdVecSize_g-1 downto 0);
       
	   i_stop_req            :in   std_logic;
	   mtime_over			 :in   std_logic;
       
       rd_en_adc_fifo_1      :in   std_logic;
       rd_en_adc_fifo_2      :in   std_logic;
       
       adc_fifo_empty_1      :out  std_logic;
       adc_fifo_empty_2      :out  std_logic;
       
       adc_fifo_data_out_1   :out std_logic_vector(11 downto 0);
       adc_fifo_data_out_2   :out std_logic_vector(11 downto 0);
       
       rd_en_peak_fifo_1     :in   std_logic;
       rd_en_peak_fifo_2     :in   std_logic;
       
       peak_fifo_empty_1     :out  std_logic;
       peak_fifo_empty_2     :out  std_logic;
       
       peak_fifo_data_out_1  :out std_logic_vector(11 downto 0);
       peak_fifo_data_out_2  :out std_logic_vector(11 downto 0)
       
         );

end entity DataCtrl;
--============================================================================
-- Entity declaration section end
--****************************************************************************


--****************************************************************************
-- Architecture definition section start - RTL
--============================================================================
architecture DataCtrl_RTL of DataCtrl is
attribute syn_noprune : boolean;
attribute syn_noprune of DataCtrl_RTL : architecture is true;
attribute syn_preserve : boolean;
attribute syn_preserve of DataCtrl_RTL: architecture is true;
  --+----------
  -- Constants, types and signals declarations start here for the architecture
  --+----------
  
  signal DATA1           :std_logic_vector(WdVecSize_g-5 downto 0);
  signal DATARDY1        :std_logic;
  signal DATA2           :std_logic_vector(WdVecSize_g-5 downto 0);
  signal DATARDY2        :std_logic;
  
  signal PEAK_FL_C1_s        :std_logic;
  signal PEAK_FL_C1_s_pos    :std_logic;
  signal PEAK_C1_s           :std_logic_vector(WdVecSize_g-5 downto 0);
  signal PEAK_C1_s_pos       :std_logic_vector(WdVecSize_g-5 downto 0);
  
  signal ADC_D1_s         :std_logic_vector(11 downto 0);
  signal ADC_DR1_s        :std_logic;
               
  signal ADC_D2_s         :std_logic_vector(11 downto 0);   
  signal ADC_DR2_s        :std_logic;

  signal i_reset_n        :std_logic;
  
  signal wr_en_adc_fifo_1   :std_logic;
  signal wr_en_adc_fifo_2   :std_logic;
  
  signal adc_fifo_data_in_1 :std_logic_vector(11 downto 0);
  signal adc_fifo_data_in_2 :std_logic_vector(11 downto 0);
        
  signal adc_fifo_full_1    :std_logic;
  signal adc_fifo_full_2    :std_logic;
  
  signal adc_fifo_wr_cnt_1  :std_logic_vector(14 downto 0);
  signal adc_fifo_wr_cnt_2  :std_logic_vector(14 downto 0);
  
  signal wr_en_peak_fifo_1   :std_logic;
  signal wr_en_peak_fifo_2   :std_logic;
  
  signal peak_fifo_data_in_1 :std_logic_vector(11 downto 0);
  signal peak_fifo_data_in_2 :std_logic_vector(11 downto 0);
        
  signal peak_fifo_full_1    :std_logic;
  signal peak_fifo_full_2    :std_logic;

  signal peak_fifo_wr_cnt_1  :std_logic_vector(10 downto 0);
  signal peak_fifo_wr_cnt_2  :std_logic_vector(10 downto 0);
  signal energy_bin_954      :std_logic_vector(11 downto 0);

  type   ENERGY_BIN_TYPE is array (0 to 1023) of std_logic_vector(11 downto 0);
  signal energy_bin_pos_data  : ENERGY_BIN_TYPE;
  signal energy_bin_neg_data  : ENERGY_BIN_TYPE;  
  signal energy_bin_cnt_1 :integer range 0 to 1025:= 0; 
  signal energy_bin_cnt_2 :integer range 0 to 1025:= 0; 
  signal s_energy_bin_pos_data_954 :std_logic_vector(11 downto 0);
  
component adc_data_fifo is
port(
        CLK     : in  std_logic;
        DATA    : in  std_logic_vector(15 downto 0);
        RE      : in  std_logic;
        RESET_N : in  std_logic;
        WE      : in  std_logic;
        -- Outputs
        EMPTY   : out std_logic;
        FULL    : out std_logic;
        Q       : out std_logic_vector(11 downto 0)
);
end component adc_data_fifo;

component peak_data_fifo is
port(
        CLK     : in  std_logic;
        DATA    : in  std_logic_vector(11 downto 0);
        RE      : in  std_logic;
        RESET_N : in  std_logic;
        WE      : in  std_logic;
        -- Outputs
        EMPTY   : out std_logic;
        FULL    : out std_logic;
        Q       : out std_logic_vector(11 downto 0)
);
end component peak_data_fifo;

component TB_adc_data_fifo is
port(
        CLK     : in  std_logic;
        DATA    : in  std_logic_vector(11 downto 0);
        RE      : in  std_logic;
        RESET_N : in  std_logic;
        WE      : in  std_logic;
        -- Outputs
        EMPTY   : out std_logic;
        FULL    : out std_logic;
        Q       : out std_logic_vector(11 downto 0)
);
end component TB_adc_data_fifo;
  
component TimeStampCtrl is
  --+----------
  -- Generic declarations
  --+----------
  generic(
          DataVecSize_g   :integer := 56;
          WdVecSize_g     :integer := 16;
          ByteSize_g      :integer := 8;
          NibbleSize_g    :integer := 4
      );

  --+----------
  -- Port name declarations
  --+----------
  port   (
       CLK100        :in  std_logic;
       RST           :in  std_logic;
       DATARDY1      :in  std_logic;
       DATARDY2      :in  std_logic;
       TIMESTAMP_C1  :out std_logic_vector(DataVecSize_g-WdVecSize_g-1 downto 0);
       TIMESTAMP_C2  :out std_logic_vector(DataVecSize_g-WdVecSize_g-1 downto 0)
         );

end component TimeStampCtrl;


component PeakDetector is
  --+----------
  -- Generic declarations
  --+----------
  generic(                        
        DataVecSize_g  		      :integer := 56;
        WdVecSize_g    		      :integer := 16;
        ByteSize_g     		      :integer := 8;
        NibbleSize_g   		      :integer := 4; 

		s_E1_C1_L        	 	  :std_logic_vector(11 downto 0) := x"000"; 
		s_E1_C1_H        	 	  :std_logic_vector(11 downto 0) := x"002"; 
		s_E2_C1_H        	 	  :std_logic_vector(11 downto 0) := x"004"; 
		s_E3_C1_H        	 	  :std_logic_vector(11 downto 0) := x"006"; 
		s_E4_C1_H        	 	  :std_logic_vector(11 downto 0) := x"008"; 
		s_E5_C1_H        	 	  :std_logic_vector(11 downto 0) := x"00A"; 
		s_E6_C1_H        	 	  :std_logic_vector(11 downto 0) := x"00C"; 
		s_E7_C1_H        	 	  :std_logic_vector(11 downto 0) := x"00E"; 
		s_E8_C1_H        	 	  :std_logic_vector(11 downto 0) := x"010"; 
		s_E9_C1_H        	 	  :std_logic_vector(11 downto 0) := x"012"; 
		s_E10_C1_H       	 	  :std_logic_vector(11 downto 0) := x"014"; 
		s_E11_C1_H				  :std_logic_vector(11 downto 0) := x"016"; 
		s_E12_C1_H				  :std_logic_vector(11 downto 0) := x"018"; 
		s_E13_C1_H				  :std_logic_vector(11 downto 0) := x"01A"; 
		s_E14_C1_H				  :std_logic_vector(11 downto 0) := x"01C"; 
		s_E15_C1_H				  :std_logic_vector(11 downto 0) := x"01E"; 
		s_E16_C1_H				  :std_logic_vector(11 downto 0) := x"020"; 
		s_E17_C1_H				  :std_logic_vector(11 downto 0) := x"022"; 
		s_E18_C1_H				  :std_logic_vector(11 downto 0) := x"024"; 
		s_E19_C1_H				  :std_logic_vector(11 downto 0) := x"026"; 
		s_E20_C1_H				  :std_logic_vector(11 downto 0) := x"028"; 
		s_E21_C1_H				  :std_logic_vector(11 downto 0) := x"02A"; 
		s_E22_C1_H				  :std_logic_vector(11 downto 0) := x"02C"; 
		s_E23_C1_H				  :std_logic_vector(11 downto 0) := x"02E"; 
		s_E24_C1_H				  :std_logic_vector(11 downto 0) := x"030"; 
		s_E25_C1_H				  :std_logic_vector(11 downto 0) := x"032"; 
		s_E26_C1_H				  :std_logic_vector(11 downto 0) := x"034"; 
		s_E27_C1_H				  :std_logic_vector(11 downto 0) := x"036"; 
		s_E28_C1_H				  :std_logic_vector(11 downto 0) := x"038"; 
		s_E29_C1_H				  :std_logic_vector(11 downto 0) := x"03A"; 
		s_E30_C1_H				  :std_logic_vector(11 downto 0) := x"03C"; 
		s_E31_C1_H				  :std_logic_vector(11 downto 0) := x"03E"; 
		s_E32_C1_H				  :std_logic_vector(11 downto 0) := x"040"; 
		s_E33_C1_H				  :std_logic_vector(11 downto 0) := x"042"; 
		s_E34_C1_H				  :std_logic_vector(11 downto 0) := x"044"; 
		s_E35_C1_H				  :std_logic_vector(11 downto 0) := x"046"; 
		s_E36_C1_H				  :std_logic_vector(11 downto 0) := x"048"; 
		s_E37_C1_H				  :std_logic_vector(11 downto 0) := x"04A"; 
		s_E38_C1_H				  :std_logic_vector(11 downto 0) := x"04C"; 
		s_E39_C1_H				  :std_logic_vector(11 downto 0) := x"04E"; 
		s_E40_C1_H				  :std_logic_vector(11 downto 0) := x"050"; 
		s_E41_C1_H				  :std_logic_vector(11 downto 0) := x"052"; 
		s_E42_C1_H				  :std_logic_vector(11 downto 0) := x"054"; 
		s_E43_C1_H				  :std_logic_vector(11 downto 0) := x"056"; 
		s_E44_C1_H				  :std_logic_vector(11 downto 0) := x"058"; 
		s_E45_C1_H				  :std_logic_vector(11 downto 0) := x"05A"; 
		s_E46_C1_H				  :std_logic_vector(11 downto 0) := x"05C"; 
		s_E47_C1_H				  :std_logic_vector(11 downto 0) := x"05E"; 
		s_E48_C1_H				  :std_logic_vector(11 downto 0) := x"060"; 
		s_E49_C1_H				  :std_logic_vector(11 downto 0) := x"062"; 
		s_E50_C1_H				  :std_logic_vector(11 downto 0) := x"064"; 
		s_E51_C1_H				  :std_logic_vector(11 downto 0) := x"066"; 
		s_E52_C1_H				  :std_logic_vector(11 downto 0) := x"068"; 
		s_E53_C1_H				  :std_logic_vector(11 downto 0) := x"06A"; 
		s_E54_C1_H				  :std_logic_vector(11 downto 0) := x"06C"; 
		s_E55_C1_H				  :std_logic_vector(11 downto 0) := x"06E"; 
		s_E56_C1_H				  :std_logic_vector(11 downto 0) := x"070"; 
		s_E57_C1_H				  :std_logic_vector(11 downto 0) := x"072"; 
		s_E58_C1_H				  :std_logic_vector(11 downto 0) := x"074"; 
		s_E59_C1_H				  :std_logic_vector(11 downto 0) := x"076"; 
		s_E60_C1_H				  :std_logic_vector(11 downto 0) := x"078"; 
		s_E61_C1_H				  :std_logic_vector(11 downto 0) := x"07A"; 
		s_E62_C1_H				  :std_logic_vector(11 downto 0) := x"07C"; 
		s_E63_C1_H				  :std_logic_vector(11 downto 0) := x"07E"; 
		s_E64_C1_H				  :std_logic_vector(11 downto 0) := x"080"; 
		s_E65_C1_H				  :std_logic_vector(11 downto 0) := x"082"; 
		s_E66_C1_H				  :std_logic_vector(11 downto 0) := x"084"; 
		s_E67_C1_H				  :std_logic_vector(11 downto 0) := x"086"; 
		s_E68_C1_H				  :std_logic_vector(11 downto 0) := x"088"; 
		s_E69_C1_H				  :std_logic_vector(11 downto 0) := x"08A"; 
		s_E70_C1_H				  :std_logic_vector(11 downto 0) := x"08C"; 
		s_E71_C1_H				  :std_logic_vector(11 downto 0) := x"08E"; 
		s_E72_C1_H				  :std_logic_vector(11 downto 0) := x"090"; 
		s_E73_C1_H				  :std_logic_vector(11 downto 0) := x"092"; 
		s_E74_C1_H				  :std_logic_vector(11 downto 0) := x"094"; 
		s_E75_C1_H				  :std_logic_vector(11 downto 0) := x"096"; 
		s_E76_C1_H				  :std_logic_vector(11 downto 0) := x"098"; 
		s_E77_C1_H				  :std_logic_vector(11 downto 0) := x"09A"; 
		s_E78_C1_H				  :std_logic_vector(11 downto 0) := x"09C"; 
		s_E79_C1_H				  :std_logic_vector(11 downto 0) := x"09E"; 
		s_E80_C1_H				  :std_logic_vector(11 downto 0) := x"0A0"; 
		s_E81_C1_H				  :std_logic_vector(11 downto 0) := x"0A2"; 
		s_E82_C1_H				  :std_logic_vector(11 downto 0) := x"0A4"; 
		s_E83_C1_H				  :std_logic_vector(11 downto 0) := x"0A6"; 
		s_E84_C1_H				  :std_logic_vector(11 downto 0) := x"0A8"; 
		s_E85_C1_H				  :std_logic_vector(11 downto 0) := x"0AA"; 
		s_E86_C1_H				  :std_logic_vector(11 downto 0) := x"0AC"; 
		s_E87_C1_H				  :std_logic_vector(11 downto 0) := x"0AE"; 
		s_E88_C1_H				  :std_logic_vector(11 downto 0) := x"0B0"; 
		s_E89_C1_H				  :std_logic_vector(11 downto 0) := x"0B2"; 
		s_E90_C1_H				  :std_logic_vector(11 downto 0) := x"0B4"; 
		s_E91_C1_H				  :std_logic_vector(11 downto 0) := x"0B6"; 
		s_E92_C1_H				  :std_logic_vector(11 downto 0) := x"0B8"; 
		s_E93_C1_H				  :std_logic_vector(11 downto 0) := x"0BA"; 
		s_E94_C1_H				  :std_logic_vector(11 downto 0) := x"0BC"; 
		s_E95_C1_H				  :std_logic_vector(11 downto 0) := x"0BE"; 
		s_E96_C1_H				  :std_logic_vector(11 downto 0) := x"0C0"; 
		s_E97_C1_H				  :std_logic_vector(11 downto 0) := x"0C2"; 
		s_E98_C1_H				  :std_logic_vector(11 downto 0) := x"0C4"; 
		s_E99_C1_H				  :std_logic_vector(11 downto 0) := x"0C6"; 
		s_E100_C1_H				  :std_logic_vector(11 downto 0) := x"0C8"; 
		s_E101_C1_H				  :std_logic_vector(11 downto 0) := x"0CA"; 
		s_E102_C1_H				  :std_logic_vector(11 downto 0) := x"0CC"; 
		s_E103_C1_H				  :std_logic_vector(11 downto 0) := x"0CE"; 
		s_E104_C1_H				  :std_logic_vector(11 downto 0) := x"0D0"; 
		s_E105_C1_H				  :std_logic_vector(11 downto 0) := x"0D2"; 
		s_E106_C1_H				  :std_logic_vector(11 downto 0) := x"0D4"; 
		s_E107_C1_H				  :std_logic_vector(11 downto 0) := x"0D6"; 
		s_E108_C1_H				  :std_logic_vector(11 downto 0) := x"0D8"; 
		s_E109_C1_H				  :std_logic_vector(11 downto 0) := x"0DA"; 
		s_E110_C1_H				  :std_logic_vector(11 downto 0) := x"0DC"; 
		s_E111_C1_H				  :std_logic_vector(11 downto 0) := x"0DE"; 
		s_E112_C1_H				  :std_logic_vector(11 downto 0) := x"0E0"; 
		s_E113_C1_H				  :std_logic_vector(11 downto 0) := x"0E2"; 
		s_E114_C1_H				  :std_logic_vector(11 downto 0) := x"0E4"; 
		s_E115_C1_H				  :std_logic_vector(11 downto 0) := x"0E6"; 
		s_E116_C1_H				  :std_logic_vector(11 downto 0) := x"0E8"; 
		s_E117_C1_H				  :std_logic_vector(11 downto 0) := x"0EA"; 
		s_E118_C1_H				  :std_logic_vector(11 downto 0) := x"0EC"; 
		s_E119_C1_H				  :std_logic_vector(11 downto 0) := x"0EE"; 
		s_E120_C1_H				  :std_logic_vector(11 downto 0) := x"0F0"; 
		s_E121_C1_H				  :std_logic_vector(11 downto 0) := x"0F2"; 
		s_E122_C1_H				  :std_logic_vector(11 downto 0) := x"0F4"; 
		s_E123_C1_H				  :std_logic_vector(11 downto 0) := x"0F6"; 
		s_E124_C1_H				  :std_logic_vector(11 downto 0) := x"0F8"; 
		s_E125_C1_H				  :std_logic_vector(11 downto 0) := x"0FA"; 
		s_E126_C1_H				  :std_logic_vector(11 downto 0) := x"0FC"; 
		s_E127_C1_H				  :std_logic_vector(11 downto 0) := x"0FE"; 
		s_E128_C1_H				  :std_logic_vector(11 downto 0) := x"100"; 
		s_E129_C1_H				  :std_logic_vector(11 downto 0) := x"102"; 
		s_E130_C1_H				  :std_logic_vector(11 downto 0) := x"104"; 
		s_E131_C1_H				  :std_logic_vector(11 downto 0) := x"106"; 
		s_E132_C1_H				  :std_logic_vector(11 downto 0) := x"108"; 
		s_E133_C1_H				  :std_logic_vector(11 downto 0) := x"10A"; 
		s_E134_C1_H				  :std_logic_vector(11 downto 0) := x"10C"; 
		s_E135_C1_H				  :std_logic_vector(11 downto 0) := x"10E"; 
		s_E136_C1_H				  :std_logic_vector(11 downto 0) := x"110"; 
		s_E137_C1_H				  :std_logic_vector(11 downto 0) := x"112"; 
		s_E138_C1_H				  :std_logic_vector(11 downto 0) := x"114"; 
		s_E139_C1_H				  :std_logic_vector(11 downto 0) := x"116"; 
		s_E140_C1_H				  :std_logic_vector(11 downto 0) := x"118"; 
		s_E141_C1_H				  :std_logic_vector(11 downto 0) := x"11A"; 
		s_E142_C1_H				  :std_logic_vector(11 downto 0) := x"11C"; 
		s_E143_C1_H				  :std_logic_vector(11 downto 0) := x"11E"; 
		s_E144_C1_H				  :std_logic_vector(11 downto 0) := x"120"; 
		s_E145_C1_H				  :std_logic_vector(11 downto 0) := x"122"; 
		s_E146_C1_H				  :std_logic_vector(11 downto 0) := x"124"; 
		s_E147_C1_H				  :std_logic_vector(11 downto 0) := x"126"; 
		s_E148_C1_H				  :std_logic_vector(11 downto 0) := x"128"; 
		s_E149_C1_H				  :std_logic_vector(11 downto 0) := x"12A"; 
		s_E150_C1_H				  :std_logic_vector(11 downto 0) := x"12C"; 
		s_E151_C1_H				  :std_logic_vector(11 downto 0) := x"12E"; 
		s_E152_C1_H				  :std_logic_vector(11 downto 0) := x"130"; 
		s_E153_C1_H				  :std_logic_vector(11 downto 0) := x"132"; 
		s_E154_C1_H				  :std_logic_vector(11 downto 0) := x"134"; 
		s_E155_C1_H				  :std_logic_vector(11 downto 0) := x"136"; 
		s_E156_C1_H				  :std_logic_vector(11 downto 0) := x"138"; 
		s_E157_C1_H				  :std_logic_vector(11 downto 0) := x"13A"; 
		s_E158_C1_H				  :std_logic_vector(11 downto 0) := x"13C"; 
		s_E159_C1_H				  :std_logic_vector(11 downto 0) := x"13E"; 
		s_E160_C1_H				  :std_logic_vector(11 downto 0) := x"140"; 
		s_E161_C1_H				  :std_logic_vector(11 downto 0) := x"142"; 
		s_E162_C1_H				  :std_logic_vector(11 downto 0) := x"144"; 
		s_E163_C1_H				  :std_logic_vector(11 downto 0) := x"146"; 
		s_E164_C1_H				  :std_logic_vector(11 downto 0) := x"148"; 
		s_E165_C1_H				  :std_logic_vector(11 downto 0) := x"14A"; 
		s_E166_C1_H				  :std_logic_vector(11 downto 0) := x"14C"; 
		s_E167_C1_H				  :std_logic_vector(11 downto 0) := x"14E"; 
		s_E168_C1_H				  :std_logic_vector(11 downto 0) := x"150"; 
		s_E169_C1_H				  :std_logic_vector(11 downto 0) := x"152"; 
		s_E170_C1_H				  :std_logic_vector(11 downto 0) := x"154"; 
		s_E171_C1_H				  :std_logic_vector(11 downto 0) := x"156"; 
		s_E172_C1_H				  :std_logic_vector(11 downto 0) := x"158"; 
		s_E173_C1_H				  :std_logic_vector(11 downto 0) := x"15A"; 
		s_E174_C1_H				  :std_logic_vector(11 downto 0) := x"15C"; 
		s_E175_C1_H				  :std_logic_vector(11 downto 0) := x"15E"; 
		s_E176_C1_H				  :std_logic_vector(11 downto 0) := x"160"; 
		s_E177_C1_H				  :std_logic_vector(11 downto 0) := x"162"; 
		s_E178_C1_H				  :std_logic_vector(11 downto 0) := x"164"; 
		s_E179_C1_H				  :std_logic_vector(11 downto 0) := x"166"; 
		s_E180_C1_H				  :std_logic_vector(11 downto 0) := x"168"; 
		s_E181_C1_H				  :std_logic_vector(11 downto 0) := x"16A"; 
		s_E182_C1_H				  :std_logic_vector(11 downto 0) := x"16C"; 
		s_E183_C1_H				  :std_logic_vector(11 downto 0) := x"16E"; 
		s_E184_C1_H				  :std_logic_vector(11 downto 0) := x"170"; 
		s_E185_C1_H				  :std_logic_vector(11 downto 0) := x"172"; 
		s_E186_C1_H				  :std_logic_vector(11 downto 0) := x"174"; 
		s_E187_C1_H				  :std_logic_vector(11 downto 0) := x"176"; 
		s_E188_C1_H				  :std_logic_vector(11 downto 0) := x"178"; 
		s_E189_C1_H				  :std_logic_vector(11 downto 0) := x"17A"; 
		s_E190_C1_H				  :std_logic_vector(11 downto 0) := x"17C"; 
		s_E191_C1_H				  :std_logic_vector(11 downto 0) := x"17E"; 
		s_E192_C1_H				  :std_logic_vector(11 downto 0) := x"180"; 
		s_E193_C1_H				  :std_logic_vector(11 downto 0) := x"182"; 
		s_E194_C1_H				  :std_logic_vector(11 downto 0) := x"184"; 
		s_E195_C1_H				  :std_logic_vector(11 downto 0) := x"186"; 
		s_E196_C1_H				  :std_logic_vector(11 downto 0) := x"188"; 
		s_E197_C1_H				  :std_logic_vector(11 downto 0) := x"18A"; 
		s_E198_C1_H				  :std_logic_vector(11 downto 0) := x"18C"; 
		s_E199_C1_H				  :std_logic_vector(11 downto 0) := x"18E"; 
		s_E200_C1_H				  :std_logic_vector(11 downto 0) := x"190"; 
		s_E201_C1_H				  :std_logic_vector(11 downto 0) := x"192"; 
		s_E202_C1_H				  :std_logic_vector(11 downto 0) := x"194"; 
		s_E203_C1_H				  :std_logic_vector(11 downto 0) := x"196"; 
		s_E204_C1_H				  :std_logic_vector(11 downto 0) := x"198"; 
		s_E205_C1_H				  :std_logic_vector(11 downto 0) := x"19A"; 
		s_E206_C1_H				  :std_logic_vector(11 downto 0) := x"19C"; 
		s_E207_C1_H				  :std_logic_vector(11 downto 0) := x"19E"; 
		s_E208_C1_H				  :std_logic_vector(11 downto 0) := x"1A0"; 
		s_E209_C1_H				  :std_logic_vector(11 downto 0) := x"1A2"; 
		s_E210_C1_H				  :std_logic_vector(11 downto 0) := x"1A4"; 
		s_E211_C1_H				  :std_logic_vector(11 downto 0) := x"1A6"; 
		s_E212_C1_H				  :std_logic_vector(11 downto 0) := x"1A8"; 
		s_E213_C1_H				  :std_logic_vector(11 downto 0) := x"1AA"; 
		s_E214_C1_H				  :std_logic_vector(11 downto 0) := x"1AC"; 
		s_E215_C1_H				  :std_logic_vector(11 downto 0) := x"1AE"; 
		s_E216_C1_H				  :std_logic_vector(11 downto 0) := x"1B0"; 
		s_E217_C1_H				  :std_logic_vector(11 downto 0) := x"1B2"; 
		s_E218_C1_H				  :std_logic_vector(11 downto 0) := x"1B4"; 
		s_E219_C1_H				  :std_logic_vector(11 downto 0) := x"1B6"; 
		s_E220_C1_H				  :std_logic_vector(11 downto 0) := x"1B8"; 
		s_E221_C1_H				  :std_logic_vector(11 downto 0) := x"1BA"; 
		s_E222_C1_H				  :std_logic_vector(11 downto 0) := x"1BC"; 
		s_E223_C1_H				  :std_logic_vector(11 downto 0) := x"1BE"; 
		s_E224_C1_H				  :std_logic_vector(11 downto 0) := x"1C0"; 
		s_E225_C1_H				  :std_logic_vector(11 downto 0) := x"1C2"; 
		s_E226_C1_H				  :std_logic_vector(11 downto 0) := x"1C4"; 
		s_E227_C1_H				  :std_logic_vector(11 downto 0) := x"1C6"; 
		s_E228_C1_H				  :std_logic_vector(11 downto 0) := x"1C8"; 
		s_E229_C1_H				  :std_logic_vector(11 downto 0) := x"1CA"; 
		s_E230_C1_H				  :std_logic_vector(11 downto 0) := x"1CC"; 
		s_E231_C1_H				  :std_logic_vector(11 downto 0) := x"1CE"; 
		s_E232_C1_H				  :std_logic_vector(11 downto 0) := x"1D0"; 
		s_E233_C1_H				  :std_logic_vector(11 downto 0) := x"1D2"; 
		s_E234_C1_H				  :std_logic_vector(11 downto 0) := x"1D4"; 
		s_E235_C1_H				  :std_logic_vector(11 downto 0) := x"1D6"; 
		s_E236_C1_H				  :std_logic_vector(11 downto 0) := x"1D8"; 
		s_E237_C1_H				  :std_logic_vector(11 downto 0) := x"1DA"; 
		s_E238_C1_H				  :std_logic_vector(11 downto 0) := x"1DC"; 
		s_E239_C1_H				  :std_logic_vector(11 downto 0) := x"1DE"; 
		s_E240_C1_H				  :std_logic_vector(11 downto 0) := x"1E0"; 
		s_E241_C1_H				  :std_logic_vector(11 downto 0) := x"1E2"; 
		s_E242_C1_H				  :std_logic_vector(11 downto 0) := x"1E4"; 
		s_E243_C1_H				  :std_logic_vector(11 downto 0) := x"1E6"; 
		s_E244_C1_H				  :std_logic_vector(11 downto 0) := x"1E8"; 
		s_E245_C1_H				  :std_logic_vector(11 downto 0) := x"1EA"; 
		s_E246_C1_H				  :std_logic_vector(11 downto 0) := x"1EC"; 
		s_E247_C1_H				  :std_logic_vector(11 downto 0) := x"1EE"; 
		s_E248_C1_H				  :std_logic_vector(11 downto 0) := x"1F0"; 
		s_E249_C1_H				  :std_logic_vector(11 downto 0) := x"1F2"; 
		s_E250_C1_H				  :std_logic_vector(11 downto 0) := x"1F4"; 
		s_E251_C1_H				  :std_logic_vector(11 downto 0) := x"1F6"; 
		s_E252_C1_H				  :std_logic_vector(11 downto 0) := x"1F8"; 
		s_E253_C1_H				  :std_logic_vector(11 downto 0) := x"1FA"; 
		s_E254_C1_H				  :std_logic_vector(11 downto 0) := x"1FC"; 
		s_E255_C1_H				  :std_logic_vector(11 downto 0) := x"1FE"; 
		s_E256_C1_H				  :std_logic_vector(11 downto 0) := x"200"; 
		s_E257_C1_H				  :std_logic_vector(11 downto 0) := x"202"; 
		s_E258_C1_H				  :std_logic_vector(11 downto 0) := x"204"; 
		s_E259_C1_H				  :std_logic_vector(11 downto 0) := x"206"; 
		s_E260_C1_H				  :std_logic_vector(11 downto 0) := x"208"; 
		s_E261_C1_H				  :std_logic_vector(11 downto 0) := x"20A"; 
		s_E262_C1_H				  :std_logic_vector(11 downto 0) := x"20C"; 
		s_E263_C1_H				  :std_logic_vector(11 downto 0) := x"20E"; 
		s_E264_C1_H				  :std_logic_vector(11 downto 0) := x"210"; 
		s_E265_C1_H				  :std_logic_vector(11 downto 0) := x"212"; 
		s_E266_C1_H				  :std_logic_vector(11 downto 0) := x"214"; 
		s_E267_C1_H				  :std_logic_vector(11 downto 0) := x"216"; 
		s_E268_C1_H				  :std_logic_vector(11 downto 0) := x"218"; 
		s_E269_C1_H				  :std_logic_vector(11 downto 0) := x"21A"; 
		s_E270_C1_H				  :std_logic_vector(11 downto 0) := x"21C"; 
		s_E271_C1_H				  :std_logic_vector(11 downto 0) := x"21E"; 
		s_E272_C1_H				  :std_logic_vector(11 downto 0) := x"220"; 
		s_E273_C1_H				  :std_logic_vector(11 downto 0) := x"222"; 
		s_E274_C1_H				  :std_logic_vector(11 downto 0) := x"224"; 
		s_E275_C1_H				  :std_logic_vector(11 downto 0) := x"226"; 
		s_E276_C1_H				  :std_logic_vector(11 downto 0) := x"228"; 
		s_E277_C1_H				  :std_logic_vector(11 downto 0) := x"22A"; 
		s_E278_C1_H				  :std_logic_vector(11 downto 0) := x"22C"; 
		s_E279_C1_H				  :std_logic_vector(11 downto 0) := x"22E"; 
		s_E280_C1_H				  :std_logic_vector(11 downto 0) := x"230"; 
		s_E281_C1_H				  :std_logic_vector(11 downto 0) := x"232"; 
		s_E282_C1_H				  :std_logic_vector(11 downto 0) := x"234"; 
		s_E283_C1_H				  :std_logic_vector(11 downto 0) := x"236"; 
		s_E284_C1_H				  :std_logic_vector(11 downto 0) := x"238"; 
		s_E285_C1_H				  :std_logic_vector(11 downto 0) := x"23A"; 
		s_E286_C1_H				  :std_logic_vector(11 downto 0) := x"23C"; 
		s_E287_C1_H				  :std_logic_vector(11 downto 0) := x"23E"; 
		s_E288_C1_H				  :std_logic_vector(11 downto 0) := x"240"; 
		s_E289_C1_H				  :std_logic_vector(11 downto 0) := x"242"; 
		s_E290_C1_H				  :std_logic_vector(11 downto 0) := x"244"; 
		s_E291_C1_H				  :std_logic_vector(11 downto 0) := x"246"; 
		s_E292_C1_H				  :std_logic_vector(11 downto 0) := x"248"; 
		s_E293_C1_H				  :std_logic_vector(11 downto 0) := x"24A"; 
		s_E294_C1_H				  :std_logic_vector(11 downto 0) := x"24C"; 
		s_E295_C1_H				  :std_logic_vector(11 downto 0) := x"24E"; 
		s_E296_C1_H				  :std_logic_vector(11 downto 0) := x"250"; 
		s_E297_C1_H				  :std_logic_vector(11 downto 0) := x"252"; 
		s_E298_C1_H				  :std_logic_vector(11 downto 0) := x"254"; 
		s_E299_C1_H				  :std_logic_vector(11 downto 0) := x"256"; 
		s_E300_C1_H				  :std_logic_vector(11 downto 0) := x"258"; 
		s_E301_C1_H				  :std_logic_vector(11 downto 0) := x"25A"; 
		s_E302_C1_H				  :std_logic_vector(11 downto 0) := x"25C"; 
		s_E303_C1_H				  :std_logic_vector(11 downto 0) := x"25E"; 
		s_E304_C1_H				  :std_logic_vector(11 downto 0) := x"260"; 
		s_E305_C1_H				  :std_logic_vector(11 downto 0) := x"262"; 
		s_E306_C1_H				  :std_logic_vector(11 downto 0) := x"264"; 
		s_E307_C1_H				  :std_logic_vector(11 downto 0) := x"266"; 
		s_E308_C1_H				  :std_logic_vector(11 downto 0) := x"268"; 
		s_E309_C1_H				  :std_logic_vector(11 downto 0) := x"26A"; 
		s_E310_C1_H				  :std_logic_vector(11 downto 0) := x"26C"; 
		s_E311_C1_H				  :std_logic_vector(11 downto 0) := x"26E"; 
		s_E312_C1_H				  :std_logic_vector(11 downto 0) := x"270"; 
		s_E313_C1_H				  :std_logic_vector(11 downto 0) := x"272"; 
		s_E314_C1_H				  :std_logic_vector(11 downto 0) := x"274"; 
		s_E315_C1_H				  :std_logic_vector(11 downto 0) := x"276"; 
		s_E316_C1_H				  :std_logic_vector(11 downto 0) := x"278"; 
		s_E317_C1_H				  :std_logic_vector(11 downto 0) := x"27A"; 
		s_E318_C1_H				  :std_logic_vector(11 downto 0) := x"27C"; 
		s_E319_C1_H				  :std_logic_vector(11 downto 0) := x"27E"; 
		s_E320_C1_H				  :std_logic_vector(11 downto 0) := x"280"; 
		s_E321_C1_H				  :std_logic_vector(11 downto 0) := x"282"; 
		s_E322_C1_H				  :std_logic_vector(11 downto 0) := x"284"; 
		s_E323_C1_H				  :std_logic_vector(11 downto 0) := x"286"; 
		s_E324_C1_H				  :std_logic_vector(11 downto 0) := x"288"; 
		s_E325_C1_H				  :std_logic_vector(11 downto 0) := x"28A"; 
		s_E326_C1_H				  :std_logic_vector(11 downto 0) := x"28C"; 
		s_E327_C1_H				  :std_logic_vector(11 downto 0) := x"28E"; 
		s_E328_C1_H				  :std_logic_vector(11 downto 0) := x"290"; 
		s_E329_C1_H				  :std_logic_vector(11 downto 0) := x"292"; 
		s_E330_C1_H				  :std_logic_vector(11 downto 0) := x"294"; 
		s_E331_C1_H				  :std_logic_vector(11 downto 0) := x"296"; 
		s_E332_C1_H				  :std_logic_vector(11 downto 0) := x"298"; 
		s_E333_C1_H				  :std_logic_vector(11 downto 0) := x"29A"; 
		s_E334_C1_H				  :std_logic_vector(11 downto 0) := x"29C"; 
		s_E335_C1_H				  :std_logic_vector(11 downto 0) := x"29E"; 
		s_E336_C1_H				  :std_logic_vector(11 downto 0) := x"2A0"; 
		s_E337_C1_H				  :std_logic_vector(11 downto 0) := x"2A2"; 
		s_E338_C1_H				  :std_logic_vector(11 downto 0) := x"2A4"; 
		s_E339_C1_H				  :std_logic_vector(11 downto 0) := x"2A6"; 
		s_E340_C1_H				  :std_logic_vector(11 downto 0) := x"2A8"; 
		s_E341_C1_H				  :std_logic_vector(11 downto 0) := x"2AA"; 
		s_E342_C1_H				  :std_logic_vector(11 downto 0) := x"2AC"; 
		s_E343_C1_H				  :std_logic_vector(11 downto 0) := x"2AE"; 
		s_E344_C1_H				  :std_logic_vector(11 downto 0) := x"2B0"; 
		s_E345_C1_H				  :std_logic_vector(11 downto 0) := x"2B2"; 
		s_E346_C1_H				  :std_logic_vector(11 downto 0) := x"2B4"; 
		s_E347_C1_H				  :std_logic_vector(11 downto 0) := x"2B6"; 
		s_E348_C1_H				  :std_logic_vector(11 downto 0) := x"2B8"; 
		s_E349_C1_H				  :std_logic_vector(11 downto 0) := x"2BA"; 
		s_E350_C1_H				  :std_logic_vector(11 downto 0) := x"2BC"; 
		s_E351_C1_H				  :std_logic_vector(11 downto 0) := x"2BE"; 
		s_E352_C1_H				  :std_logic_vector(11 downto 0) := x"2C0"; 
		s_E353_C1_H				  :std_logic_vector(11 downto 0) := x"2C2"; 
		s_E354_C1_H				  :std_logic_vector(11 downto 0) := x"2C4"; 
		s_E355_C1_H				  :std_logic_vector(11 downto 0) := x"2C6"; 
		s_E356_C1_H				  :std_logic_vector(11 downto 0) := x"2C8"; 
		s_E357_C1_H				  :std_logic_vector(11 downto 0) := x"2CA"; 
		s_E358_C1_H				  :std_logic_vector(11 downto 0) := x"2CC"; 
		s_E359_C1_H				  :std_logic_vector(11 downto 0) := x"2CE"; 
		s_E360_C1_H				  :std_logic_vector(11 downto 0) := x"2D0"; 
		s_E361_C1_H				  :std_logic_vector(11 downto 0) := x"2D2"; 
		s_E362_C1_H				  :std_logic_vector(11 downto 0) := x"2D4"; 
		s_E363_C1_H				  :std_logic_vector(11 downto 0) := x"2D6"; 
		s_E364_C1_H				  :std_logic_vector(11 downto 0) := x"2D8"; 
		s_E365_C1_H				  :std_logic_vector(11 downto 0) := x"2DA"; 
		s_E366_C1_H				  :std_logic_vector(11 downto 0) := x"2DC"; 
		s_E367_C1_H				  :std_logic_vector(11 downto 0) := x"2DE"; 
		s_E368_C1_H				  :std_logic_vector(11 downto 0) := x"2E0"; 
		s_E369_C1_H				  :std_logic_vector(11 downto 0) := x"2E2"; 
		s_E370_C1_H				  :std_logic_vector(11 downto 0) := x"2E4"; 
		s_E371_C1_H				  :std_logic_vector(11 downto 0) := x"2E6"; 
		s_E372_C1_H				  :std_logic_vector(11 downto 0) := x"2E8"; 
		s_E373_C1_H				  :std_logic_vector(11 downto 0) := x"2EA"; 
		s_E374_C1_H				  :std_logic_vector(11 downto 0) := x"2EC"; 
		s_E375_C1_H				  :std_logic_vector(11 downto 0) := x"2EE"; 
		s_E376_C1_H				  :std_logic_vector(11 downto 0) := x"2F0"; 
		s_E377_C1_H				  :std_logic_vector(11 downto 0) := x"2F2"; 
		s_E378_C1_H				  :std_logic_vector(11 downto 0) := x"2F4"; 
		s_E379_C1_H				  :std_logic_vector(11 downto 0) := x"2F6"; 
		s_E380_C1_H				  :std_logic_vector(11 downto 0) := x"2F8"; 
		s_E381_C1_H				  :std_logic_vector(11 downto 0) := x"2FA"; 
		s_E382_C1_H				  :std_logic_vector(11 downto 0) := x"2FC"; 
		s_E383_C1_H				  :std_logic_vector(11 downto 0) := x"2FE"; 
		s_E384_C1_H				  :std_logic_vector(11 downto 0) := x"300"; 
		s_E385_C1_H				  :std_logic_vector(11 downto 0) := x"302"; 
		s_E386_C1_H				  :std_logic_vector(11 downto 0) := x"304"; 
		s_E387_C1_H				  :std_logic_vector(11 downto 0) := x"306"; 
		s_E388_C1_H				  :std_logic_vector(11 downto 0) := x"308"; 
		s_E389_C1_H				  :std_logic_vector(11 downto 0) := x"30A"; 
		s_E390_C1_H				  :std_logic_vector(11 downto 0) := x"30C"; 
		s_E391_C1_H				  :std_logic_vector(11 downto 0) := x"30E"; 
		s_E392_C1_H				  :std_logic_vector(11 downto 0) := x"310"; 
		s_E393_C1_H				  :std_logic_vector(11 downto 0) := x"312"; 
		s_E394_C1_H				  :std_logic_vector(11 downto 0) := x"314"; 
		s_E395_C1_H				  :std_logic_vector(11 downto 0) := x"316"; 
		s_E396_C1_H				  :std_logic_vector(11 downto 0) := x"318"; 
		s_E397_C1_H				  :std_logic_vector(11 downto 0) := x"31A"; 
		s_E398_C1_H				  :std_logic_vector(11 downto 0) := x"31C"; 
		s_E399_C1_H				  :std_logic_vector(11 downto 0) := x"31E"; 
		s_E400_C1_H				  :std_logic_vector(11 downto 0) := x"320"; 
		s_E401_C1_H				  :std_logic_vector(11 downto 0) := x"322"; 
		s_E402_C1_H				  :std_logic_vector(11 downto 0) := x"324"; 
		s_E403_C1_H				  :std_logic_vector(11 downto 0) := x"326"; 
		s_E404_C1_H				  :std_logic_vector(11 downto 0) := x"328"; 
		s_E405_C1_H				  :std_logic_vector(11 downto 0) := x"32A"; 
		s_E406_C1_H				  :std_logic_vector(11 downto 0) := x"32C"; 
		s_E407_C1_H				  :std_logic_vector(11 downto 0) := x"32E"; 
		s_E408_C1_H				  :std_logic_vector(11 downto 0) := x"330"; 
		s_E409_C1_H				  :std_logic_vector(11 downto 0) := x"332"; 
		s_E410_C1_H				  :std_logic_vector(11 downto 0) := x"334"; 
		s_E411_C1_H				  :std_logic_vector(11 downto 0) := x"336"; 
		s_E412_C1_H				  :std_logic_vector(11 downto 0) := x"338"; 
		s_E413_C1_H				  :std_logic_vector(11 downto 0) := x"33A"; 
		s_E414_C1_H				  :std_logic_vector(11 downto 0) := x"33C"; 
		s_E415_C1_H				  :std_logic_vector(11 downto 0) := x"33E"; 
		s_E416_C1_H				  :std_logic_vector(11 downto 0) := x"340"; 
		s_E417_C1_H				  :std_logic_vector(11 downto 0) := x"342"; 
		s_E418_C1_H				  :std_logic_vector(11 downto 0) := x"344"; 
		s_E419_C1_H				  :std_logic_vector(11 downto 0) := x"346"; 
		s_E420_C1_H				  :std_logic_vector(11 downto 0) := x"348"; 
		s_E421_C1_H				  :std_logic_vector(11 downto 0) := x"34A"; 
		s_E422_C1_H				  :std_logic_vector(11 downto 0) := x"34C"; 
		s_E423_C1_H				  :std_logic_vector(11 downto 0) := x"34E"; 
		s_E424_C1_H				  :std_logic_vector(11 downto 0) := x"350"; 
		s_E425_C1_H				  :std_logic_vector(11 downto 0) := x"352"; 
		s_E426_C1_H				  :std_logic_vector(11 downto 0) := x"354"; 
		s_E427_C1_H				  :std_logic_vector(11 downto 0) := x"356"; 
		s_E428_C1_H				  :std_logic_vector(11 downto 0) := x"358"; 
		s_E429_C1_H				  :std_logic_vector(11 downto 0) := x"35A"; 
		s_E430_C1_H				  :std_logic_vector(11 downto 0) := x"35C"; 
		s_E431_C1_H				  :std_logic_vector(11 downto 0) := x"35E"; 
		s_E432_C1_H				  :std_logic_vector(11 downto 0) := x"360"; 
		s_E433_C1_H				  :std_logic_vector(11 downto 0) := x"362"; 
		s_E434_C1_H				  :std_logic_vector(11 downto 0) := x"364"; 
		s_E435_C1_H				  :std_logic_vector(11 downto 0) := x"366"; 
		s_E436_C1_H				  :std_logic_vector(11 downto 0) := x"368"; 
		s_E437_C1_H				  :std_logic_vector(11 downto 0) := x"36A"; 
		s_E438_C1_H				  :std_logic_vector(11 downto 0) := x"36C"; 
		s_E439_C1_H				  :std_logic_vector(11 downto 0) := x"36E"; 
		s_E440_C1_H				  :std_logic_vector(11 downto 0) := x"370"; 
		s_E441_C1_H				  :std_logic_vector(11 downto 0) := x"372"; 
		s_E442_C1_H				  :std_logic_vector(11 downto 0) := x"374"; 
		s_E443_C1_H				  :std_logic_vector(11 downto 0) := x"376"; 
		s_E444_C1_H				  :std_logic_vector(11 downto 0) := x"378"; 
		s_E445_C1_H				  :std_logic_vector(11 downto 0) := x"37A"; 
		s_E446_C1_H				  :std_logic_vector(11 downto 0) := x"37C"; 
		s_E447_C1_H				  :std_logic_vector(11 downto 0) := x"37E"; 
		s_E448_C1_H				  :std_logic_vector(11 downto 0) := x"380"; 
		s_E449_C1_H				  :std_logic_vector(11 downto 0) := x"382"; 
		s_E450_C1_H				  :std_logic_vector(11 downto 0) := x"384"; 
		s_E451_C1_H				  :std_logic_vector(11 downto 0) := x"386"; 
		s_E452_C1_H				  :std_logic_vector(11 downto 0) := x"388"; 
		s_E453_C1_H				  :std_logic_vector(11 downto 0) := x"38A"; 
		s_E454_C1_H				  :std_logic_vector(11 downto 0) := x"38C"; 
		s_E455_C1_H				  :std_logic_vector(11 downto 0) := x"38E"; 
		s_E456_C1_H				  :std_logic_vector(11 downto 0) := x"390"; 
		s_E457_C1_H				  :std_logic_vector(11 downto 0) := x"392"; 
		s_E458_C1_H				  :std_logic_vector(11 downto 0) := x"394"; 
		s_E459_C1_H				  :std_logic_vector(11 downto 0) := x"396"; 
		s_E460_C1_H				  :std_logic_vector(11 downto 0) := x"398"; 
		s_E461_C1_H				  :std_logic_vector(11 downto 0) := x"39A"; 
		s_E462_C1_H				  :std_logic_vector(11 downto 0) := x"39C"; 
		s_E463_C1_H				  :std_logic_vector(11 downto 0) := x"39E"; 
		s_E464_C1_H				  :std_logic_vector(11 downto 0) := x"3A0"; 
		s_E465_C1_H				  :std_logic_vector(11 downto 0) := x"3A2"; 
		s_E466_C1_H				  :std_logic_vector(11 downto 0) := x"3A4"; 
		s_E467_C1_H				  :std_logic_vector(11 downto 0) := x"3A6"; 
		s_E468_C1_H				  :std_logic_vector(11 downto 0) := x"3A8"; 
		s_E469_C1_H				  :std_logic_vector(11 downto 0) := x"3AA"; 
		s_E470_C1_H				  :std_logic_vector(11 downto 0) := x"3AC"; 
		s_E471_C1_H				  :std_logic_vector(11 downto 0) := x"3AE"; 
		s_E472_C1_H				  :std_logic_vector(11 downto 0) := x"3B0"; 
		s_E473_C1_H				  :std_logic_vector(11 downto 0) := x"3B2"; 
		s_E474_C1_H				  :std_logic_vector(11 downto 0) := x"3B4"; 
		s_E475_C1_H				  :std_logic_vector(11 downto 0) := x"3B6"; 
		s_E476_C1_H				  :std_logic_vector(11 downto 0) := x"3B8"; 
		s_E477_C1_H				  :std_logic_vector(11 downto 0) := x"3BA"; 
		s_E478_C1_H				  :std_logic_vector(11 downto 0) := x"3BC"; 
		s_E479_C1_H				  :std_logic_vector(11 downto 0) := x"3BE"; 
		s_E480_C1_H				  :std_logic_vector(11 downto 0) := x"3C0"; 
		s_E481_C1_H				  :std_logic_vector(11 downto 0) := x"3C2"; 
		s_E482_C1_H				  :std_logic_vector(11 downto 0) := x"3C4"; 
		s_E483_C1_H				  :std_logic_vector(11 downto 0) := x"3C6"; 
		s_E484_C1_H				  :std_logic_vector(11 downto 0) := x"3C8"; 
		s_E485_C1_H				  :std_logic_vector(11 downto 0) := x"3CA"; 
		s_E486_C1_H				  :std_logic_vector(11 downto 0) := x"3CC"; 
		s_E487_C1_H				  :std_logic_vector(11 downto 0) := x"3CE"; 
		s_E488_C1_H				  :std_logic_vector(11 downto 0) := x"3D0"; 
		s_E489_C1_H				  :std_logic_vector(11 downto 0) := x"3D2"; 
		s_E490_C1_H				  :std_logic_vector(11 downto 0) := x"3D4"; 
		s_E491_C1_H				  :std_logic_vector(11 downto 0) := x"3D6"; 
		s_E492_C1_H				  :std_logic_vector(11 downto 0) := x"3D8"; 
		s_E493_C1_H				  :std_logic_vector(11 downto 0) := x"3DA"; 
		s_E494_C1_H				  :std_logic_vector(11 downto 0) := x"3DC"; 
		s_E495_C1_H				  :std_logic_vector(11 downto 0) := x"3DE"; 
		s_E496_C1_H				  :std_logic_vector(11 downto 0) := x"3E0"; 
		s_E497_C1_H				  :std_logic_vector(11 downto 0) := x"3E2"; 
		s_E498_C1_H				  :std_logic_vector(11 downto 0) := x"3E4"; 
		s_E499_C1_H				  :std_logic_vector(11 downto 0) := x"3E6"; 
		s_E500_C1_H				  :std_logic_vector(11 downto 0) := x"3E8"; 
		s_E501_C1_H				  :std_logic_vector(11 downto 0) := x"3EA"; 
		s_E502_C1_H				  :std_logic_vector(11 downto 0) := x"3EC"; 
		s_E503_C1_H				  :std_logic_vector(11 downto 0) := x"3EE"; 
		s_E504_C1_H				  :std_logic_vector(11 downto 0) := x"3F0"; 
		s_E505_C1_H				  :std_logic_vector(11 downto 0) := x"3F2"; 
		s_E506_C1_H				  :std_logic_vector(11 downto 0) := x"3F4"; 
		s_E507_C1_H				  :std_logic_vector(11 downto 0) := x"3F6"; 
		s_E508_C1_H				  :std_logic_vector(11 downto 0) := x"3F8"; 
		s_E509_C1_H				  :std_logic_vector(11 downto 0) := x"3FA"; 
		s_E510_C1_H				  :std_logic_vector(11 downto 0) := x"3FC"; 
		s_E511_C1_H				  :std_logic_vector(11 downto 0) := x"3FE"; 
		s_E512_C1_H				  :std_logic_vector(11 downto 0) := x"400"; 
		s_E513_C1_H				  :std_logic_vector(11 downto 0) := x"402"; 
		s_E514_C1_H				  :std_logic_vector(11 downto 0) := x"404"; 
		s_E515_C1_H				  :std_logic_vector(11 downto 0) := x"406"; 
		s_E516_C1_H				  :std_logic_vector(11 downto 0) := x"408"; 
		s_E517_C1_H				  :std_logic_vector(11 downto 0) := x"40A"; 
		s_E518_C1_H				  :std_logic_vector(11 downto 0) := x"40C"; 
		s_E519_C1_H				  :std_logic_vector(11 downto 0) := x"40E"; 
		s_E520_C1_H				  :std_logic_vector(11 downto 0) := x"410"; 
		s_E521_C1_H				  :std_logic_vector(11 downto 0) := x"412"; 
		s_E522_C1_H				  :std_logic_vector(11 downto 0) := x"414"; 
		s_E523_C1_H				  :std_logic_vector(11 downto 0) := x"416"; 
		s_E524_C1_H				  :std_logic_vector(11 downto 0) := x"418"; 
		s_E525_C1_H				  :std_logic_vector(11 downto 0) := x"41A"; 
		s_E526_C1_H				  :std_logic_vector(11 downto 0) := x"41C"; 
		s_E527_C1_H				  :std_logic_vector(11 downto 0) := x"41E"; 
		s_E528_C1_H				  :std_logic_vector(11 downto 0) := x"420"; 
		s_E529_C1_H				  :std_logic_vector(11 downto 0) := x"422"; 
		s_E530_C1_H				  :std_logic_vector(11 downto 0) := x"424"; 
		s_E531_C1_H				  :std_logic_vector(11 downto 0) := x"426"; 
		s_E532_C1_H				  :std_logic_vector(11 downto 0) := x"428"; 
		s_E533_C1_H				  :std_logic_vector(11 downto 0) := x"42A"; 
		s_E534_C1_H				  :std_logic_vector(11 downto 0) := x"42C"; 
		s_E535_C1_H				  :std_logic_vector(11 downto 0) := x"42E"; 
		s_E536_C1_H				  :std_logic_vector(11 downto 0) := x"430"; 
		s_E537_C1_H				  :std_logic_vector(11 downto 0) := x"432"; 
		s_E538_C1_H				  :std_logic_vector(11 downto 0) := x"434"; 
		s_E539_C1_H				  :std_logic_vector(11 downto 0) := x"436"; 
		s_E540_C1_H				  :std_logic_vector(11 downto 0) := x"438"; 
		s_E541_C1_H				  :std_logic_vector(11 downto 0) := x"43A"; 
		s_E542_C1_H				  :std_logic_vector(11 downto 0) := x"43C"; 
		s_E543_C1_H				  :std_logic_vector(11 downto 0) := x"43E"; 
		s_E544_C1_H				  :std_logic_vector(11 downto 0) := x"440"; 
		s_E545_C1_H				  :std_logic_vector(11 downto 0) := x"442"; 
		s_E546_C1_H				  :std_logic_vector(11 downto 0) := x"444"; 
		s_E547_C1_H				  :std_logic_vector(11 downto 0) := x"446"; 
		s_E548_C1_H				  :std_logic_vector(11 downto 0) := x"448"; 
		s_E549_C1_H				  :std_logic_vector(11 downto 0) := x"44A"; 
		s_E550_C1_H				  :std_logic_vector(11 downto 0) := x"44C"; 
		s_E551_C1_H				  :std_logic_vector(11 downto 0) := x"44E"; 
		s_E552_C1_H				  :std_logic_vector(11 downto 0) := x"450"; 
		s_E553_C1_H				  :std_logic_vector(11 downto 0) := x"452"; 
		s_E554_C1_H				  :std_logic_vector(11 downto 0) := x"454"; 
		s_E555_C1_H				  :std_logic_vector(11 downto 0) := x"456"; 
		s_E556_C1_H				  :std_logic_vector(11 downto 0) := x"458"; 
		s_E557_C1_H				  :std_logic_vector(11 downto 0) := x"45A"; 
		s_E558_C1_H				  :std_logic_vector(11 downto 0) := x"45C"; 
		s_E559_C1_H				  :std_logic_vector(11 downto 0) := x"45E"; 
		s_E560_C1_H				  :std_logic_vector(11 downto 0) := x"460"; 
		s_E561_C1_H				  :std_logic_vector(11 downto 0) := x"462"; 
		s_E562_C1_H				  :std_logic_vector(11 downto 0) := x"464"; 
		s_E563_C1_H				  :std_logic_vector(11 downto 0) := x"466"; 
		s_E564_C1_H				  :std_logic_vector(11 downto 0) := x"468"; 
		s_E565_C1_H				  :std_logic_vector(11 downto 0) := x"46A"; 
		s_E566_C1_H				  :std_logic_vector(11 downto 0) := x"46C"; 
		s_E567_C1_H				  :std_logic_vector(11 downto 0) := x"46E"; 
		s_E568_C1_H				  :std_logic_vector(11 downto 0) := x"470"; 
		s_E569_C1_H				  :std_logic_vector(11 downto 0) := x"472"; 
		s_E570_C1_H				  :std_logic_vector(11 downto 0) := x"474"; 
		s_E571_C1_H				  :std_logic_vector(11 downto 0) := x"476"; 
		s_E572_C1_H				  :std_logic_vector(11 downto 0) := x"478"; 
		s_E573_C1_H				  :std_logic_vector(11 downto 0) := x"47A"; 
		s_E574_C1_H				  :std_logic_vector(11 downto 0) := x"47C"; 
		s_E575_C1_H				  :std_logic_vector(11 downto 0) := x"47E"; 
		s_E576_C1_H				  :std_logic_vector(11 downto 0) := x"480"; 
		s_E577_C1_H				  :std_logic_vector(11 downto 0) := x"482"; 
		s_E578_C1_H				  :std_logic_vector(11 downto 0) := x"484"; 
		s_E579_C1_H				  :std_logic_vector(11 downto 0) := x"486"; 
		s_E580_C1_H				  :std_logic_vector(11 downto 0) := x"488"; 
		s_E581_C1_H				  :std_logic_vector(11 downto 0) := x"48A"; 
		s_E582_C1_H				  :std_logic_vector(11 downto 0) := x"48C"; 
		s_E583_C1_H				  :std_logic_vector(11 downto 0) := x"48E"; 
		s_E584_C1_H				  :std_logic_vector(11 downto 0) := x"490"; 
		s_E585_C1_H				  :std_logic_vector(11 downto 0) := x"492"; 
		s_E586_C1_H				  :std_logic_vector(11 downto 0) := x"494"; 
		s_E587_C1_H				  :std_logic_vector(11 downto 0) := x"496"; 
		s_E588_C1_H				  :std_logic_vector(11 downto 0) := x"498"; 
		s_E589_C1_H				  :std_logic_vector(11 downto 0) := x"49A"; 
		s_E590_C1_H				  :std_logic_vector(11 downto 0) := x"49C"; 
		s_E591_C1_H				  :std_logic_vector(11 downto 0) := x"49E"; 
		s_E592_C1_H				  :std_logic_vector(11 downto 0) := x"4A0"; 
		s_E593_C1_H				  :std_logic_vector(11 downto 0) := x"4A2"; 
		s_E594_C1_H				  :std_logic_vector(11 downto 0) := x"4A4"; 
		s_E595_C1_H				  :std_logic_vector(11 downto 0) := x"4A6"; 
		s_E596_C1_H				  :std_logic_vector(11 downto 0) := x"4A8"; 
		s_E597_C1_H				  :std_logic_vector(11 downto 0) := x"4AA"; 
		s_E598_C1_H				  :std_logic_vector(11 downto 0) := x"4AC"; 
		s_E599_C1_H				  :std_logic_vector(11 downto 0) := x"4AE"; 
		s_E600_C1_H				  :std_logic_vector(11 downto 0) := x"4B0"; 
		s_E601_C1_H				  :std_logic_vector(11 downto 0) := x"4B2"; 
		s_E602_C1_H				  :std_logic_vector(11 downto 0) := x"4B4"; 
		s_E603_C1_H				  :std_logic_vector(11 downto 0) := x"4B6"; 
		s_E604_C1_H				  :std_logic_vector(11 downto 0) := x"4B8"; 
		s_E605_C1_H				  :std_logic_vector(11 downto 0) := x"4BA"; 
		s_E606_C1_H				  :std_logic_vector(11 downto 0) := x"4BC"; 
		s_E607_C1_H				  :std_logic_vector(11 downto 0) := x"4BE"; 
		s_E608_C1_H				  :std_logic_vector(11 downto 0) := x"4C0"; 
		s_E609_C1_H				  :std_logic_vector(11 downto 0) := x"4C2"; 
		s_E610_C1_H				  :std_logic_vector(11 downto 0) := x"4C4"; 
		s_E611_C1_H				  :std_logic_vector(11 downto 0) := x"4C6"; 
		s_E612_C1_H				  :std_logic_vector(11 downto 0) := x"4C8"; 
		s_E613_C1_H				  :std_logic_vector(11 downto 0) := x"4CA"; 
		s_E614_C1_H				  :std_logic_vector(11 downto 0) := x"4CC"; 
		s_E615_C1_H				  :std_logic_vector(11 downto 0) := x"4CE"; 
		s_E616_C1_H				  :std_logic_vector(11 downto 0) := x"4D0"; 
		s_E617_C1_H				  :std_logic_vector(11 downto 0) := x"4D2"; 
		s_E618_C1_H				  :std_logic_vector(11 downto 0) := x"4D4"; 
		s_E619_C1_H				  :std_logic_vector(11 downto 0) := x"4D6"; 
		s_E620_C1_H				  :std_logic_vector(11 downto 0) := x"4D8"; 
		s_E621_C1_H				  :std_logic_vector(11 downto 0) := x"4DA"; 
		s_E622_C1_H				  :std_logic_vector(11 downto 0) := x"4DC"; 
		s_E623_C1_H				  :std_logic_vector(11 downto 0) := x"4DE"; 
		s_E624_C1_H				  :std_logic_vector(11 downto 0) := x"4E0"; 
		s_E625_C1_H				  :std_logic_vector(11 downto 0) := x"4E2"; 
		s_E626_C1_H				  :std_logic_vector(11 downto 0) := x"4E4"; 
		s_E627_C1_H				  :std_logic_vector(11 downto 0) := x"4E6"; 
		s_E628_C1_H				  :std_logic_vector(11 downto 0) := x"4E8"; 
		s_E629_C1_H				  :std_logic_vector(11 downto 0) := x"4EA"; 
		s_E630_C1_H				  :std_logic_vector(11 downto 0) := x"4EC"; 
		s_E631_C1_H				  :std_logic_vector(11 downto 0) := x"4EE"; 
		s_E632_C1_H				  :std_logic_vector(11 downto 0) := x"4F0"; 
		s_E633_C1_H				  :std_logic_vector(11 downto 0) := x"4F2"; 
		s_E634_C1_H				  :std_logic_vector(11 downto 0) := x"4F4"; 
		s_E635_C1_H				  :std_logic_vector(11 downto 0) := x"4F6"; 
		s_E636_C1_H				  :std_logic_vector(11 downto 0) := x"4F8"; 
		s_E637_C1_H				  :std_logic_vector(11 downto 0) := x"4FA"; 
		s_E638_C1_H				  :std_logic_vector(11 downto 0) := x"4FC"; 
		s_E639_C1_H				  :std_logic_vector(11 downto 0) := x"4FE"; 
		s_E640_C1_H				  :std_logic_vector(11 downto 0) := x"500"; 
		s_E641_C1_H				  :std_logic_vector(11 downto 0) := x"502"; 
		s_E642_C1_H				  :std_logic_vector(11 downto 0) := x"504"; 
		s_E643_C1_H				  :std_logic_vector(11 downto 0) := x"506"; 
		s_E644_C1_H				  :std_logic_vector(11 downto 0) := x"508"; 
		s_E645_C1_H				  :std_logic_vector(11 downto 0) := x"50A"; 
		s_E646_C1_H				  :std_logic_vector(11 downto 0) := x"50C"; 
		s_E647_C1_H				  :std_logic_vector(11 downto 0) := x"50E"; 
		s_E648_C1_H				  :std_logic_vector(11 downto 0) := x"510"; 
		s_E649_C1_H				  :std_logic_vector(11 downto 0) := x"512"; 
		s_E650_C1_H				  :std_logic_vector(11 downto 0) := x"514"; 
		s_E651_C1_H				  :std_logic_vector(11 downto 0) := x"516"; 
		s_E652_C1_H				  :std_logic_vector(11 downto 0) := x"518"; 
		s_E653_C1_H				  :std_logic_vector(11 downto 0) := x"51A"; 
		s_E654_C1_H				  :std_logic_vector(11 downto 0) := x"51C"; 
		s_E655_C1_H				  :std_logic_vector(11 downto 0) := x"51E"; 
		s_E656_C1_H				  :std_logic_vector(11 downto 0) := x"520"; 
		s_E657_C1_H				  :std_logic_vector(11 downto 0) := x"522"; 
		s_E658_C1_H				  :std_logic_vector(11 downto 0) := x"524"; 
		s_E659_C1_H				  :std_logic_vector(11 downto 0) := x"526"; 
		s_E660_C1_H				  :std_logic_vector(11 downto 0) := x"528"; 
		s_E661_C1_H				  :std_logic_vector(11 downto 0) := x"52A"; 
		s_E662_C1_H				  :std_logic_vector(11 downto 0) := x"52C"; 
		s_E663_C1_H				  :std_logic_vector(11 downto 0) := x"52E"; 
		s_E664_C1_H				  :std_logic_vector(11 downto 0) := x"530"; 
		s_E665_C1_H				  :std_logic_vector(11 downto 0) := x"532"; 
		s_E666_C1_H				  :std_logic_vector(11 downto 0) := x"534"; 
		s_E667_C1_H				  :std_logic_vector(11 downto 0) := x"536"; 
		s_E668_C1_H				  :std_logic_vector(11 downto 0) := x"538"; 
		s_E669_C1_H				  :std_logic_vector(11 downto 0) := x"53A"; 
		s_E670_C1_H				  :std_logic_vector(11 downto 0) := x"53C"; 
		s_E671_C1_H				  :std_logic_vector(11 downto 0) := x"53E"; 
		s_E672_C1_H				  :std_logic_vector(11 downto 0) := x"540"; 
		s_E673_C1_H				  :std_logic_vector(11 downto 0) := x"542"; 
		s_E674_C1_H				  :std_logic_vector(11 downto 0) := x"544"; 
		s_E675_C1_H				  :std_logic_vector(11 downto 0) := x"546"; 
		s_E676_C1_H				  :std_logic_vector(11 downto 0) := x"548"; 
		s_E677_C1_H				  :std_logic_vector(11 downto 0) := x"54A"; 
		s_E678_C1_H				  :std_logic_vector(11 downto 0) := x"54C"; 
		s_E679_C1_H				  :std_logic_vector(11 downto 0) := x"54E"; 
		s_E680_C1_H				  :std_logic_vector(11 downto 0) := x"550"; 
		s_E681_C1_H				  :std_logic_vector(11 downto 0) := x"552"; 
		s_E682_C1_H				  :std_logic_vector(11 downto 0) := x"554"; 
		s_E683_C1_H				  :std_logic_vector(11 downto 0) := x"556"; 
		s_E684_C1_H				  :std_logic_vector(11 downto 0) := x"558"; 
		s_E685_C1_H				  :std_logic_vector(11 downto 0) := x"55A"; 
		s_E686_C1_H				  :std_logic_vector(11 downto 0) := x"55C"; 
		s_E687_C1_H				  :std_logic_vector(11 downto 0) := x"55E"; 
		s_E688_C1_H				  :std_logic_vector(11 downto 0) := x"560"; 
		s_E689_C1_H				  :std_logic_vector(11 downto 0) := x"562"; 
		s_E690_C1_H				  :std_logic_vector(11 downto 0) := x"564"; 
		s_E691_C1_H				  :std_logic_vector(11 downto 0) := x"566"; 
		s_E692_C1_H				  :std_logic_vector(11 downto 0) := x"568"; 
		s_E693_C1_H				  :std_logic_vector(11 downto 0) := x"56A"; 
		s_E694_C1_H				  :std_logic_vector(11 downto 0) := x"56C"; 
		s_E695_C1_H				  :std_logic_vector(11 downto 0) := x"56E"; 
		s_E696_C1_H				  :std_logic_vector(11 downto 0) := x"570"; 
		s_E697_C1_H				  :std_logic_vector(11 downto 0) := x"572"; 
		s_E698_C1_H				  :std_logic_vector(11 downto 0) := x"574"; 
		s_E699_C1_H				  :std_logic_vector(11 downto 0) := x"576"; 
		s_E700_C1_H				  :std_logic_vector(11 downto 0) := x"578"; 
		s_E701_C1_H				  :std_logic_vector(11 downto 0) := x"57A"; 
		s_E702_C1_H				  :std_logic_vector(11 downto 0) := x"57C"; 
		s_E703_C1_H				  :std_logic_vector(11 downto 0) := x"57E"; 
		s_E704_C1_H				  :std_logic_vector(11 downto 0) := x"580"; 
		s_E705_C1_H				  :std_logic_vector(11 downto 0) := x"582"; 
		s_E706_C1_H				  :std_logic_vector(11 downto 0) := x"584"; 
		s_E707_C1_H				  :std_logic_vector(11 downto 0) := x"586"; 
		s_E708_C1_H				  :std_logic_vector(11 downto 0) := x"588"; 
		s_E709_C1_H				  :std_logic_vector(11 downto 0) := x"58A"; 
		s_E710_C1_H				  :std_logic_vector(11 downto 0) := x"58C"; 
		s_E711_C1_H				  :std_logic_vector(11 downto 0) := x"58E"; 
		s_E712_C1_H				  :std_logic_vector(11 downto 0) := x"590"; 
		s_E713_C1_H				  :std_logic_vector(11 downto 0) := x"592"; 
		s_E714_C1_H				  :std_logic_vector(11 downto 0) := x"594"; 
		s_E715_C1_H				  :std_logic_vector(11 downto 0) := x"596"; 
		s_E716_C1_H				  :std_logic_vector(11 downto 0) := x"598"; 
		s_E717_C1_H				  :std_logic_vector(11 downto 0) := x"59A"; 
		s_E718_C1_H				  :std_logic_vector(11 downto 0) := x"59C"; 
		s_E719_C1_H				  :std_logic_vector(11 downto 0) := x"59E"; 
		s_E720_C1_H				  :std_logic_vector(11 downto 0) := x"5A0"; 
		s_E721_C1_H				  :std_logic_vector(11 downto 0) := x"5A2"; 
		s_E722_C1_H				  :std_logic_vector(11 downto 0) := x"5A4"; 
		s_E723_C1_H				  :std_logic_vector(11 downto 0) := x"5A6"; 
		s_E724_C1_H				  :std_logic_vector(11 downto 0) := x"5A8"; 
		s_E725_C1_H				  :std_logic_vector(11 downto 0) := x"5AA"; 
		s_E726_C1_H				  :std_logic_vector(11 downto 0) := x"5AC"; 
		s_E727_C1_H				  :std_logic_vector(11 downto 0) := x"5AE"; 
		s_E728_C1_H				  :std_logic_vector(11 downto 0) := x"5B0"; 
		s_E729_C1_H				  :std_logic_vector(11 downto 0) := x"5B2"; 
		s_E730_C1_H				  :std_logic_vector(11 downto 0) := x"5B4"; 
		s_E731_C1_H				  :std_logic_vector(11 downto 0) := x"5B6"; 
		s_E732_C1_H				  :std_logic_vector(11 downto 0) := x"5B8"; 
		s_E733_C1_H				  :std_logic_vector(11 downto 0) := x"5BA"; 
		s_E734_C1_H				  :std_logic_vector(11 downto 0) := x"5BC"; 
		s_E735_C1_H				  :std_logic_vector(11 downto 0) := x"5BE"; 
		s_E736_C1_H				  :std_logic_vector(11 downto 0) := x"5C0"; 
		s_E737_C1_H				  :std_logic_vector(11 downto 0) := x"5C2"; 
		s_E738_C1_H				  :std_logic_vector(11 downto 0) := x"5C4"; 
		s_E739_C1_H				  :std_logic_vector(11 downto 0) := x"5C6"; 
		s_E740_C1_H				  :std_logic_vector(11 downto 0) := x"5C8"; 
		s_E741_C1_H				  :std_logic_vector(11 downto 0) := x"5CA"; 
		s_E742_C1_H				  :std_logic_vector(11 downto 0) := x"5CC"; 
		s_E743_C1_H				  :std_logic_vector(11 downto 0) := x"5CE"; 
		s_E744_C1_H				  :std_logic_vector(11 downto 0) := x"5D0"; 
		s_E745_C1_H				  :std_logic_vector(11 downto 0) := x"5D2"; 
		s_E746_C1_H				  :std_logic_vector(11 downto 0) := x"5D4"; 
		s_E747_C1_H				  :std_logic_vector(11 downto 0) := x"5D6"; 
		s_E748_C1_H				  :std_logic_vector(11 downto 0) := x"5D8"; 
		s_E749_C1_H				  :std_logic_vector(11 downto 0) := x"5DA"; 
		s_E750_C1_H				  :std_logic_vector(11 downto 0) := x"5DC"; 
		s_E751_C1_H				  :std_logic_vector(11 downto 0) := x"5DE"; 
		s_E752_C1_H				  :std_logic_vector(11 downto 0) := x"5E0"; 
		s_E753_C1_H				  :std_logic_vector(11 downto 0) := x"5E2"; 
		s_E754_C1_H				  :std_logic_vector(11 downto 0) := x"5E4"; 
		s_E755_C1_H				  :std_logic_vector(11 downto 0) := x"5E6"; 
		s_E756_C1_H				  :std_logic_vector(11 downto 0) := x"5E8"; 
		s_E757_C1_H				  :std_logic_vector(11 downto 0) := x"5EA"; 
		s_E758_C1_H				  :std_logic_vector(11 downto 0) := x"5EC"; 
		s_E759_C1_H				  :std_logic_vector(11 downto 0) := x"5EE"; 
		s_E760_C1_H				  :std_logic_vector(11 downto 0) := x"5F0"; 
		s_E761_C1_H				  :std_logic_vector(11 downto 0) := x"5F2"; 
		s_E762_C1_H				  :std_logic_vector(11 downto 0) := x"5F4"; 
		s_E763_C1_H				  :std_logic_vector(11 downto 0) := x"5F6"; 
		s_E764_C1_H				  :std_logic_vector(11 downto 0) := x"5F8"; 
		s_E765_C1_H				  :std_logic_vector(11 downto 0) := x"5FA"; 
		s_E766_C1_H				  :std_logic_vector(11 downto 0) := x"5FC"; 
		s_E767_C1_H				  :std_logic_vector(11 downto 0) := x"5FE"; 
		s_E768_C1_H				  :std_logic_vector(11 downto 0) := x"600"; 
		s_E769_C1_H				  :std_logic_vector(11 downto 0) := x"602"; 
		s_E770_C1_H				  :std_logic_vector(11 downto 0) := x"604"; 
		s_E771_C1_H				  :std_logic_vector(11 downto 0) := x"606"; 
		s_E772_C1_H				  :std_logic_vector(11 downto 0) := x"608"; 
		s_E773_C1_H				  :std_logic_vector(11 downto 0) := x"60A"; 
		s_E774_C1_H				  :std_logic_vector(11 downto 0) := x"60C"; 
		s_E775_C1_H				  :std_logic_vector(11 downto 0) := x"60E"; 
		s_E776_C1_H				  :std_logic_vector(11 downto 0) := x"610"; 
		s_E777_C1_H				  :std_logic_vector(11 downto 0) := x"612"; 
		s_E778_C1_H				  :std_logic_vector(11 downto 0) := x"614"; 
		s_E779_C1_H				  :std_logic_vector(11 downto 0) := x"616"; 
		s_E780_C1_H				  :std_logic_vector(11 downto 0) := x"618"; 
		s_E781_C1_H				  :std_logic_vector(11 downto 0) := x"61A"; 
		s_E782_C1_H				  :std_logic_vector(11 downto 0) := x"61C"; 
		s_E783_C1_H				  :std_logic_vector(11 downto 0) := x"61E"; 
		s_E784_C1_H				  :std_logic_vector(11 downto 0) := x"620"; 
		s_E785_C1_H				  :std_logic_vector(11 downto 0) := x"622"; 
		s_E786_C1_H				  :std_logic_vector(11 downto 0) := x"624"; 
		s_E787_C1_H				  :std_logic_vector(11 downto 0) := x"626"; 
		s_E788_C1_H				  :std_logic_vector(11 downto 0) := x"628"; 
		s_E789_C1_H				  :std_logic_vector(11 downto 0) := x"62A"; 
		s_E790_C1_H				  :std_logic_vector(11 downto 0) := x"62C"; 
		s_E791_C1_H				  :std_logic_vector(11 downto 0) := x"62E"; 
		s_E792_C1_H				  :std_logic_vector(11 downto 0) := x"630"; 
		s_E793_C1_H				  :std_logic_vector(11 downto 0) := x"632"; 
		s_E794_C1_H				  :std_logic_vector(11 downto 0) := x"634"; 
		s_E795_C1_H				  :std_logic_vector(11 downto 0) := x"636"; 
		s_E796_C1_H				  :std_logic_vector(11 downto 0) := x"638"; 
		s_E797_C1_H				  :std_logic_vector(11 downto 0) := x"63A"; 
		s_E798_C1_H				  :std_logic_vector(11 downto 0) := x"63C"; 
		s_E799_C1_H				  :std_logic_vector(11 downto 0) := x"63E"; 
		s_E800_C1_H				  :std_logic_vector(11 downto 0) := x"640"; 
		s_E801_C1_H				  :std_logic_vector(11 downto 0) := x"642"; 
		s_E802_C1_H				  :std_logic_vector(11 downto 0) := x"644"; 
		s_E803_C1_H				  :std_logic_vector(11 downto 0) := x"646"; 
		s_E804_C1_H				  :std_logic_vector(11 downto 0) := x"648"; 
		s_E805_C1_H				  :std_logic_vector(11 downto 0) := x"64A"; 
		s_E806_C1_H				  :std_logic_vector(11 downto 0) := x"64C"; 
		s_E807_C1_H				  :std_logic_vector(11 downto 0) := x"64E"; 
		s_E808_C1_H				  :std_logic_vector(11 downto 0) := x"650"; 
		s_E809_C1_H				  :std_logic_vector(11 downto 0) := x"652"; 
		s_E810_C1_H				  :std_logic_vector(11 downto 0) := x"654"; 
		s_E811_C1_H				  :std_logic_vector(11 downto 0) := x"656"; 
		s_E812_C1_H				  :std_logic_vector(11 downto 0) := x"658"; 
		s_E813_C1_H				  :std_logic_vector(11 downto 0) := x"65A"; 
		s_E814_C1_H				  :std_logic_vector(11 downto 0) := x"65C"; 
		s_E815_C1_H				  :std_logic_vector(11 downto 0) := x"65E"; 
		s_E816_C1_H				  :std_logic_vector(11 downto 0) := x"660"; 
		s_E817_C1_H				  :std_logic_vector(11 downto 0) := x"662"; 
		s_E818_C1_H				  :std_logic_vector(11 downto 0) := x"664"; 
		s_E819_C1_H				  :std_logic_vector(11 downto 0) := x"666"; 
		s_E820_C1_H				  :std_logic_vector(11 downto 0) := x"668"; 
		s_E821_C1_H				  :std_logic_vector(11 downto 0) := x"66A"; 
		s_E822_C1_H				  :std_logic_vector(11 downto 0) := x"66C"; 
		s_E823_C1_H				  :std_logic_vector(11 downto 0) := x"66E"; 
		s_E824_C1_H				  :std_logic_vector(11 downto 0) := x"670"; 
		s_E825_C1_H				  :std_logic_vector(11 downto 0) := x"672"; 
		s_E826_C1_H				  :std_logic_vector(11 downto 0) := x"674"; 
		s_E827_C1_H				  :std_logic_vector(11 downto 0) := x"676"; 
		s_E828_C1_H				  :std_logic_vector(11 downto 0) := x"678"; 
		s_E829_C1_H				  :std_logic_vector(11 downto 0) := x"67A"; 
		s_E830_C1_H				  :std_logic_vector(11 downto 0) := x"67C"; 
		s_E831_C1_H				  :std_logic_vector(11 downto 0) := x"67E"; 
		s_E832_C1_H				  :std_logic_vector(11 downto 0) := x"680"; 
		s_E833_C1_H				  :std_logic_vector(11 downto 0) := x"682"; 
		s_E834_C1_H				  :std_logic_vector(11 downto 0) := x"684"; 
		s_E835_C1_H				  :std_logic_vector(11 downto 0) := x"686"; 
		s_E836_C1_H				  :std_logic_vector(11 downto 0) := x"688"; 
		s_E837_C1_H				  :std_logic_vector(11 downto 0) := x"68A"; 
		s_E838_C1_H				  :std_logic_vector(11 downto 0) := x"68C"; 
		s_E839_C1_H				  :std_logic_vector(11 downto 0) := x"68E"; 
		s_E840_C1_H				  :std_logic_vector(11 downto 0) := x"690"; 
		s_E841_C1_H				  :std_logic_vector(11 downto 0) := x"692"; 
		s_E842_C1_H				  :std_logic_vector(11 downto 0) := x"694"; 
		s_E843_C1_H				  :std_logic_vector(11 downto 0) := x"696"; 
		s_E844_C1_H				  :std_logic_vector(11 downto 0) := x"698"; 
		s_E845_C1_H				  :std_logic_vector(11 downto 0) := x"69A"; 
		s_E846_C1_H				  :std_logic_vector(11 downto 0) := x"69C"; 
		s_E847_C1_H				  :std_logic_vector(11 downto 0) := x"69E"; 
		s_E848_C1_H				  :std_logic_vector(11 downto 0) := x"6A0"; 
		s_E849_C1_H				  :std_logic_vector(11 downto 0) := x"6A2"; 
		s_E850_C1_H				  :std_logic_vector(11 downto 0) := x"6A4"; 
		s_E851_C1_H				  :std_logic_vector(11 downto 0) := x"6A6"; 
		s_E852_C1_H				  :std_logic_vector(11 downto 0) := x"6A8"; 
		s_E853_C1_H				  :std_logic_vector(11 downto 0) := x"6AA"; 
		s_E854_C1_H				  :std_logic_vector(11 downto 0) := x"6AC"; 
		s_E855_C1_H				  :std_logic_vector(11 downto 0) := x"6AE"; 
		s_E856_C1_H				  :std_logic_vector(11 downto 0) := x"6B0"; 
		s_E857_C1_H				  :std_logic_vector(11 downto 0) := x"6B2"; 
		s_E858_C1_H				  :std_logic_vector(11 downto 0) := x"6B4"; 
		s_E859_C1_H				  :std_logic_vector(11 downto 0) := x"6B6"; 
		s_E860_C1_H				  :std_logic_vector(11 downto 0) := x"6B8"; 
		s_E861_C1_H				  :std_logic_vector(11 downto 0) := x"6BA"; 
		s_E862_C1_H				  :std_logic_vector(11 downto 0) := x"6BC"; 
		s_E863_C1_H				  :std_logic_vector(11 downto 0) := x"6BE"; 
		s_E864_C1_H				  :std_logic_vector(11 downto 0) := x"6C0"; 
		s_E865_C1_H				  :std_logic_vector(11 downto 0) := x"6C2"; 
		s_E866_C1_H				  :std_logic_vector(11 downto 0) := x"6C4"; 
		s_E867_C1_H				  :std_logic_vector(11 downto 0) := x"6C6"; 
		s_E868_C1_H				  :std_logic_vector(11 downto 0) := x"6C8"; 
		s_E869_C1_H				  :std_logic_vector(11 downto 0) := x"6CA"; 
		s_E870_C1_H				  :std_logic_vector(11 downto 0) := x"6CC"; 
		s_E871_C1_H				  :std_logic_vector(11 downto 0) := x"6CE"; 
		s_E872_C1_H				  :std_logic_vector(11 downto 0) := x"6D0"; 
		s_E873_C1_H				  :std_logic_vector(11 downto 0) := x"6D2"; 
		s_E874_C1_H				  :std_logic_vector(11 downto 0) := x"6D4"; 
		s_E875_C1_H				  :std_logic_vector(11 downto 0) := x"6D6"; 
		s_E876_C1_H				  :std_logic_vector(11 downto 0) := x"6D8"; 
		s_E877_C1_H				  :std_logic_vector(11 downto 0) := x"6DA"; 
		s_E878_C1_H				  :std_logic_vector(11 downto 0) := x"6DC"; 
		s_E879_C1_H				  :std_logic_vector(11 downto 0) := x"6DE"; 
		s_E880_C1_H				  :std_logic_vector(11 downto 0) := x"6E0"; 
		s_E881_C1_H				  :std_logic_vector(11 downto 0) := x"6E2"; 
		s_E882_C1_H				  :std_logic_vector(11 downto 0) := x"6E4"; 
		s_E883_C1_H				  :std_logic_vector(11 downto 0) := x"6E6"; 
		s_E884_C1_H				  :std_logic_vector(11 downto 0) := x"6E8"; 
		s_E885_C1_H				  :std_logic_vector(11 downto 0) := x"6EA"; 
		s_E886_C1_H				  :std_logic_vector(11 downto 0) := x"6EC"; 
		s_E887_C1_H				  :std_logic_vector(11 downto 0) := x"6EE"; 
		s_E888_C1_H				  :std_logic_vector(11 downto 0) := x"6F0"; 
		s_E889_C1_H				  :std_logic_vector(11 downto 0) := x"6F2"; 
		s_E890_C1_H				  :std_logic_vector(11 downto 0) := x"6F4"; 
		s_E891_C1_H				  :std_logic_vector(11 downto 0) := x"6F6"; 
		s_E892_C1_H				  :std_logic_vector(11 downto 0) := x"6F8"; 
		s_E893_C1_H				  :std_logic_vector(11 downto 0) := x"6FA"; 
		s_E894_C1_H				  :std_logic_vector(11 downto 0) := x"6FC"; 
		s_E895_C1_H				  :std_logic_vector(11 downto 0) := x"6FE"; 
		s_E896_C1_H				  :std_logic_vector(11 downto 0) := x"700"; 
		s_E897_C1_H				  :std_logic_vector(11 downto 0) := x"702"; 
		s_E898_C1_H				  :std_logic_vector(11 downto 0) := x"704"; 
		s_E899_C1_H				  :std_logic_vector(11 downto 0) := x"706"; 
		s_E900_C1_H				  :std_logic_vector(11 downto 0) := x"708"; 
		s_E901_C1_H				  :std_logic_vector(11 downto 0) := x"70A"; 
		s_E902_C1_H				  :std_logic_vector(11 downto 0) := x"70C"; 
		s_E903_C1_H				  :std_logic_vector(11 downto 0) := x"70E"; 
		s_E904_C1_H				  :std_logic_vector(11 downto 0) := x"710"; 
		s_E905_C1_H				  :std_logic_vector(11 downto 0) := x"712"; 
		s_E906_C1_H				  :std_logic_vector(11 downto 0) := x"714"; 
		s_E907_C1_H				  :std_logic_vector(11 downto 0) := x"716"; 
		s_E908_C1_H				  :std_logic_vector(11 downto 0) := x"718"; 
		s_E909_C1_H				  :std_logic_vector(11 downto 0) := x"71A"; 
		s_E910_C1_H				  :std_logic_vector(11 downto 0) := x"71C"; 
		s_E911_C1_H				  :std_logic_vector(11 downto 0) := x"71E"; 
		s_E912_C1_H				  :std_logic_vector(11 downto 0) := x"720"; 
		s_E913_C1_H				  :std_logic_vector(11 downto 0) := x"722"; 
		s_E914_C1_H				  :std_logic_vector(11 downto 0) := x"724"; 
		s_E915_C1_H				  :std_logic_vector(11 downto 0) := x"726"; 
		s_E916_C1_H				  :std_logic_vector(11 downto 0) := x"728"; 
		s_E917_C1_H				  :std_logic_vector(11 downto 0) := x"72A"; 
		s_E918_C1_H				  :std_logic_vector(11 downto 0) := x"72C"; 
		s_E919_C1_H				  :std_logic_vector(11 downto 0) := x"72E"; 
		s_E920_C1_H				  :std_logic_vector(11 downto 0) := x"730"; 
		s_E921_C1_H				  :std_logic_vector(11 downto 0) := x"732"; 
		s_E922_C1_H				  :std_logic_vector(11 downto 0) := x"734"; 
		s_E923_C1_H				  :std_logic_vector(11 downto 0) := x"736"; 
		s_E924_C1_H				  :std_logic_vector(11 downto 0) := x"738"; 
		s_E925_C1_H				  :std_logic_vector(11 downto 0) := x"73A"; 
		s_E926_C1_H				  :std_logic_vector(11 downto 0) := x"73C"; 
		s_E927_C1_H				  :std_logic_vector(11 downto 0) := x"73E"; 
		s_E928_C1_H				  :std_logic_vector(11 downto 0) := x"740"; 
		s_E929_C1_H				  :std_logic_vector(11 downto 0) := x"742"; 
		s_E930_C1_H				  :std_logic_vector(11 downto 0) := x"744"; 
		s_E931_C1_H				  :std_logic_vector(11 downto 0) := x"746"; 
		s_E932_C1_H				  :std_logic_vector(11 downto 0) := x"748"; 
		s_E933_C1_H				  :std_logic_vector(11 downto 0) := x"74A"; 
		s_E934_C1_H				  :std_logic_vector(11 downto 0) := x"74C"; 
		s_E935_C1_H				  :std_logic_vector(11 downto 0) := x"74E"; 
		s_E936_C1_H				  :std_logic_vector(11 downto 0) := x"750"; 
		s_E937_C1_H				  :std_logic_vector(11 downto 0) := x"752"; 
		s_E938_C1_H				  :std_logic_vector(11 downto 0) := x"754"; 
		s_E939_C1_H				  :std_logic_vector(11 downto 0) := x"756"; 
		s_E940_C1_H				  :std_logic_vector(11 downto 0) := x"758"; 
		s_E941_C1_H				  :std_logic_vector(11 downto 0) := x"75A"; 
		s_E942_C1_H				  :std_logic_vector(11 downto 0) := x"75C"; 
		s_E943_C1_H				  :std_logic_vector(11 downto 0) := x"75E"; 
		s_E944_C1_H				  :std_logic_vector(11 downto 0) := x"760"; 
		s_E945_C1_H				  :std_logic_vector(11 downto 0) := x"762"; 
		s_E946_C1_H				  :std_logic_vector(11 downto 0) := x"764"; 
		s_E947_C1_H				  :std_logic_vector(11 downto 0) := x"766"; 
		s_E948_C1_H				  :std_logic_vector(11 downto 0) := x"768"; 
		s_E949_C1_H				  :std_logic_vector(11 downto 0) := x"76A"; 
		s_E950_C1_H				  :std_logic_vector(11 downto 0) := x"76C"; 
		s_E951_C1_H				  :std_logic_vector(11 downto 0) := x"76E"; 
		s_E952_C1_H				  :std_logic_vector(11 downto 0) := x"770"; 
		s_E953_C1_H				  :std_logic_vector(11 downto 0) := x"772"; 
		s_E954_C1_H				  :std_logic_vector(11 downto 0) := x"774"; 
		s_E955_C1_H				  :std_logic_vector(11 downto 0) := x"776"; 
		s_E956_C1_H				  :std_logic_vector(11 downto 0) := x"778"; 
		s_E957_C1_H				  :std_logic_vector(11 downto 0) := x"77A"; 
		s_E958_C1_H				  :std_logic_vector(11 downto 0) := x"77C"; 
		s_E959_C1_H				  :std_logic_vector(11 downto 0) := x"77E"; 
		s_E960_C1_H				  :std_logic_vector(11 downto 0) := x"780"; 
		s_E961_C1_H				  :std_logic_vector(11 downto 0) := x"782"; 
		s_E962_C1_H				  :std_logic_vector(11 downto 0) := x"784"; 
		s_E963_C1_H				  :std_logic_vector(11 downto 0) := x"786"; 
		s_E964_C1_H				  :std_logic_vector(11 downto 0) := x"788"; 
		s_E965_C1_H				  :std_logic_vector(11 downto 0) := x"78A"; 
		s_E966_C1_H				  :std_logic_vector(11 downto 0) := x"78C"; 
		s_E967_C1_H				  :std_logic_vector(11 downto 0) := x"78E"; 
		s_E968_C1_H				  :std_logic_vector(11 downto 0) := x"790"; 
		s_E969_C1_H				  :std_logic_vector(11 downto 0) := x"792"; 
		s_E970_C1_H				  :std_logic_vector(11 downto 0) := x"794"; 
		s_E971_C1_H				  :std_logic_vector(11 downto 0) := x"796"; 
		s_E972_C1_H				  :std_logic_vector(11 downto 0) := x"798"; 
		s_E973_C1_H				  :std_logic_vector(11 downto 0) := x"79A"; 
		s_E974_C1_H				  :std_logic_vector(11 downto 0) := x"79C"; 
		s_E975_C1_H				  :std_logic_vector(11 downto 0) := x"79E"; 
		s_E976_C1_H				  :std_logic_vector(11 downto 0) := x"7A0"; 
		s_E977_C1_H				  :std_logic_vector(11 downto 0) := x"7A2"; 
		s_E978_C1_H				  :std_logic_vector(11 downto 0) := x"7A4"; 
		s_E979_C1_H				  :std_logic_vector(11 downto 0) := x"7A6"; 
		s_E980_C1_H				  :std_logic_vector(11 downto 0) := x"7A8"; 
		s_E981_C1_H				  :std_logic_vector(11 downto 0) := x"7AA"; 
		s_E982_C1_H				  :std_logic_vector(11 downto 0) := x"7AC"; 
		s_E983_C1_H				  :std_logic_vector(11 downto 0) := x"7AE"; 
		s_E984_C1_H				  :std_logic_vector(11 downto 0) := x"7B0"; 
		s_E985_C1_H				  :std_logic_vector(11 downto 0) := x"7B2"; 
		s_E986_C1_H				  :std_logic_vector(11 downto 0) := x"7B4"; 
		s_E987_C1_H				  :std_logic_vector(11 downto 0) := x"7B6"; 
		s_E988_C1_H				  :std_logic_vector(11 downto 0) := x"7B8"; 
		s_E989_C1_H				  :std_logic_vector(11 downto 0) := x"7BA"; 
		s_E990_C1_H				  :std_logic_vector(11 downto 0) := x"7BC"; 
		s_E991_C1_H				  :std_logic_vector(11 downto 0) := x"7BE"; 
		s_E992_C1_H				  :std_logic_vector(11 downto 0) := x"7C0"; 
		s_E993_C1_H				  :std_logic_vector(11 downto 0) := x"7C2"; 
		s_E994_C1_H				  :std_logic_vector(11 downto 0) := x"7C4"; 
		s_E995_C1_H				  :std_logic_vector(11 downto 0) := x"7C6"; 
		s_E996_C1_H				  :std_logic_vector(11 downto 0) := x"7C8"; 
		s_E997_C1_H				  :std_logic_vector(11 downto 0) := x"7CA"; 
		s_E998_C1_H				  :std_logic_vector(11 downto 0) := x"7CC"; 
		s_E999_C1_H				  :std_logic_vector(11 downto 0) := x"7CE"; 
		s_E1000_C1_H			  :std_logic_vector(11 downto 0) := x"7D0"; 
		s_E1001_C1_H			  :std_logic_vector(11 downto 0) := x"7D2"; 
		s_E1002_C1_H			  :std_logic_vector(11 downto 0) := x"7D4"; 
		s_E1003_C1_H			  :std_logic_vector(11 downto 0) := x"7D6"; 
		s_E1004_C1_H			  :std_logic_vector(11 downto 0) := x"7D8"; 
		s_E1005_C1_H			  :std_logic_vector(11 downto 0) := x"7DA"; 
		s_E1006_C1_H			  :std_logic_vector(11 downto 0) := x"7DC"; 
		s_E1007_C1_H			  :std_logic_vector(11 downto 0) := x"7DE"; 
		s_E1008_C1_H			  :std_logic_vector(11 downto 0) := x"7E0"; 
		s_E1009_C1_H			  :std_logic_vector(11 downto 0) := x"7E2"; 
		s_E1010_C1_H			  :std_logic_vector(11 downto 0) := x"7E4"; 
		s_E1011_C1_H			  :std_logic_vector(11 downto 0) := x"7E6"; 
		s_E1012_C1_H			  :std_logic_vector(11 downto 0) := x"7E8"; 
		s_E1013_C1_H			  :std_logic_vector(11 downto 0) := x"7EA"; 
		s_E1014_C1_H			  :std_logic_vector(11 downto 0) := x"7EC"; 
		s_E1015_C1_H			  :std_logic_vector(11 downto 0) := x"7EE"; 
		s_E1016_C1_H			  :std_logic_vector(11 downto 0) := x"7F0"; 
		s_E1017_C1_H			  :std_logic_vector(11 downto 0) := x"7F2"; 
		s_E1018_C1_H			  :std_logic_vector(11 downto 0) := x"7F4"; 
		s_E1019_C1_H			  :std_logic_vector(11 downto 0) := x"7F6"; 
		s_E1020_C1_H			  :std_logic_vector(11 downto 0) := x"7F8"; 
		s_E1021_C1_H			  :std_logic_vector(11 downto 0) := x"7FA"; 
		s_E1022_C1_H			  :std_logic_vector(11 downto 0) := x"7FC"; 
		s_E1023_C1_H			  :std_logic_vector(11 downto 0) := x"7FE"; 
		s_E1024_C1_H			  :std_logic_vector(11 downto 0) := x"7FF"; 
		
		s_E2_C1_L       	 	  :std_logic_vector(11 downto 0) := x"002"; 
		s_E3_C1_L       	 	  :std_logic_vector(11 downto 0) := x"004"; 
		s_E4_C1_L       	 	  :std_logic_vector(11 downto 0) := x"006"; 
		s_E5_C1_L       	 	  :std_logic_vector(11 downto 0) := x"008"; 
		s_E6_C1_L       	 	  :std_logic_vector(11 downto 0) := x"00A"; 
		s_E7_C1_L       	 	  :std_logic_vector(11 downto 0) := x"00C"; 
		s_E8_C1_L       	 	  :std_logic_vector(11 downto 0) := x"00E"; 
		s_E9_C1_L       	 	  :std_logic_vector(11 downto 0) := x"010"; 
		s_E10_C1_L       	 	  :std_logic_vector(11 downto 0) := x"012"; 
		s_E11_C1_L				  :std_logic_vector(11 downto 0) := x"014"; 
		s_E12_C1_L				  :std_logic_vector(11 downto 0) := x"016"; 
		s_E13_C1_L				  :std_logic_vector(11 downto 0) := x"018"; 
		s_E14_C1_L				  :std_logic_vector(11 downto 0) := x"01A"; 
		s_E15_C1_L				  :std_logic_vector(11 downto 0) := x"01C"; 
		s_E16_C1_L				  :std_logic_vector(11 downto 0) := x"01E"; 
		s_E17_C1_L				  :std_logic_vector(11 downto 0) := x"020"; 
		s_E18_C1_L				  :std_logic_vector(11 downto 0) := x"022"; 
		s_E19_C1_L				  :std_logic_vector(11 downto 0) := x"024"; 
		s_E20_C1_L				  :std_logic_vector(11 downto 0) := x"026"; 
		s_E21_C1_L				  :std_logic_vector(11 downto 0) := x"028"; 
		s_E22_C1_L				  :std_logic_vector(11 downto 0) := x"02A"; 
		s_E23_C1_L				  :std_logic_vector(11 downto 0) := x"02C"; 
		s_E24_C1_L				  :std_logic_vector(11 downto 0) := x"02E"; 
		s_E25_C1_L				  :std_logic_vector(11 downto 0) := x"030"; 
		s_E26_C1_L				  :std_logic_vector(11 downto 0) := x"032"; 
		s_E27_C1_L				  :std_logic_vector(11 downto 0) := x"034"; 
		s_E28_C1_L				  :std_logic_vector(11 downto 0) := x"036"; 
		s_E29_C1_L				  :std_logic_vector(11 downto 0) := x"038"; 
		s_E30_C1_L				  :std_logic_vector(11 downto 0) := x"03A"; 
		s_E31_C1_L				  :std_logic_vector(11 downto 0) := x"03C"; 
		s_E32_C1_L				  :std_logic_vector(11 downto 0) := x"03E"; 
		s_E33_C1_L				  :std_logic_vector(11 downto 0) := x"040"; 
		s_E34_C1_L				  :std_logic_vector(11 downto 0) := x"042"; 
		s_E35_C1_L				  :std_logic_vector(11 downto 0) := x"044"; 
		s_E36_C1_L				  :std_logic_vector(11 downto 0) := x"046"; 
		s_E37_C1_L				  :std_logic_vector(11 downto 0) := x"048"; 
		s_E38_C1_L				  :std_logic_vector(11 downto 0) := x"04A"; 
		s_E39_C1_L				  :std_logic_vector(11 downto 0) := x"04C"; 
		s_E40_C1_L				  :std_logic_vector(11 downto 0) := x"04E"; 
		s_E41_C1_L				  :std_logic_vector(11 downto 0) := x"050"; 
		s_E42_C1_L				  :std_logic_vector(11 downto 0) := x"052"; 
		s_E43_C1_L				  :std_logic_vector(11 downto 0) := x"054"; 
		s_E44_C1_L				  :std_logic_vector(11 downto 0) := x"056"; 
		s_E45_C1_L				  :std_logic_vector(11 downto 0) := x"058"; 
		s_E46_C1_L				  :std_logic_vector(11 downto 0) := x"05A"; 
		s_E47_C1_L				  :std_logic_vector(11 downto 0) := x"05C"; 
		s_E48_C1_L				  :std_logic_vector(11 downto 0) := x"05E"; 
		s_E49_C1_L				  :std_logic_vector(11 downto 0) := x"060"; 
		s_E50_C1_L				  :std_logic_vector(11 downto 0) := x"062"; 
		s_E51_C1_L				  :std_logic_vector(11 downto 0) := x"064"; 
		s_E52_C1_L				  :std_logic_vector(11 downto 0) := x"066"; 
		s_E53_C1_L				  :std_logic_vector(11 downto 0) := x"068"; 
		s_E54_C1_L				  :std_logic_vector(11 downto 0) := x"06A"; 
		s_E55_C1_L				  :std_logic_vector(11 downto 0) := x"06C"; 
		s_E56_C1_L				  :std_logic_vector(11 downto 0) := x"06E"; 
		s_E57_C1_L				  :std_logic_vector(11 downto 0) := x"070"; 
		s_E58_C1_L				  :std_logic_vector(11 downto 0) := x"072"; 
		s_E59_C1_L				  :std_logic_vector(11 downto 0) := x"074"; 
		s_E60_C1_L				  :std_logic_vector(11 downto 0) := x"076"; 
		s_E61_C1_L				  :std_logic_vector(11 downto 0) := x"078"; 
		s_E62_C1_L				  :std_logic_vector(11 downto 0) := x"07A"; 
		s_E63_C1_L				  :std_logic_vector(11 downto 0) := x"07C"; 
		s_E64_C1_L				  :std_logic_vector(11 downto 0) := x"07E"; 
		s_E65_C1_L				  :std_logic_vector(11 downto 0) := x"080"; 
		s_E66_C1_L				  :std_logic_vector(11 downto 0) := x"082"; 
		s_E67_C1_L				  :std_logic_vector(11 downto 0) := x"084"; 
		s_E68_C1_L				  :std_logic_vector(11 downto 0) := x"086"; 
		s_E69_C1_L				  :std_logic_vector(11 downto 0) := x"088"; 
		s_E70_C1_L				  :std_logic_vector(11 downto 0) := x"08A"; 
		s_E71_C1_L				  :std_logic_vector(11 downto 0) := x"08C"; 
		s_E72_C1_L				  :std_logic_vector(11 downto 0) := x"08E"; 
		s_E73_C1_L				  :std_logic_vector(11 downto 0) := x"090"; 
		s_E74_C1_L				  :std_logic_vector(11 downto 0) := x"092"; 
		s_E75_C1_L				  :std_logic_vector(11 downto 0) := x"094"; 
		s_E76_C1_L				  :std_logic_vector(11 downto 0) := x"096"; 
		s_E77_C1_L				  :std_logic_vector(11 downto 0) := x"098"; 
		s_E78_C1_L				  :std_logic_vector(11 downto 0) := x"09A"; 
		s_E79_C1_L				  :std_logic_vector(11 downto 0) := x"09C"; 
		s_E80_C1_L				  :std_logic_vector(11 downto 0) := x"09E"; 
		s_E81_C1_L				  :std_logic_vector(11 downto 0) := x"0A0"; 
		s_E82_C1_L				  :std_logic_vector(11 downto 0) := x"0A2"; 
		s_E83_C1_L				  :std_logic_vector(11 downto 0) := x"0A4"; 
		s_E84_C1_L				  :std_logic_vector(11 downto 0) := x"0A6"; 
		s_E85_C1_L				  :std_logic_vector(11 downto 0) := x"0A8"; 
		s_E86_C1_L				  :std_logic_vector(11 downto 0) := x"0AA"; 
		s_E87_C1_L				  :std_logic_vector(11 downto 0) := x"0AC"; 
		s_E88_C1_L				  :std_logic_vector(11 downto 0) := x"0AE"; 
		s_E89_C1_L				  :std_logic_vector(11 downto 0) := x"0B0"; 
		s_E90_C1_L				  :std_logic_vector(11 downto 0) := x"0B2"; 
		s_E91_C1_L				  :std_logic_vector(11 downto 0) := x"0B4"; 
		s_E92_C1_L				  :std_logic_vector(11 downto 0) := x"0B6"; 
		s_E93_C1_L				  :std_logic_vector(11 downto 0) := x"0B8"; 
		s_E94_C1_L				  :std_logic_vector(11 downto 0) := x"0BA"; 
		s_E95_C1_L				  :std_logic_vector(11 downto 0) := x"0BC"; 
		s_E96_C1_L				  :std_logic_vector(11 downto 0) := x"0BE"; 
		s_E97_C1_L				  :std_logic_vector(11 downto 0) := x"0C0"; 
		s_E98_C1_L				  :std_logic_vector(11 downto 0) := x"0C2"; 
		s_E99_C1_L				  :std_logic_vector(11 downto 0) := x"0C4"; 
		s_E100_C1_L				  :std_logic_vector(11 downto 0) := x"0C6"; 
		s_E101_C1_L				  :std_logic_vector(11 downto 0) := x"0C8"; 
		s_E102_C1_L				  :std_logic_vector(11 downto 0) := x"0CA"; 
		s_E103_C1_L				  :std_logic_vector(11 downto 0) := x"0CC"; 
		s_E104_C1_L				  :std_logic_vector(11 downto 0) := x"0CE"; 
		s_E105_C1_L				  :std_logic_vector(11 downto 0) := x"0D0"; 
		s_E106_C1_L				  :std_logic_vector(11 downto 0) := x"0D2"; 
		s_E107_C1_L				  :std_logic_vector(11 downto 0) := x"0D4"; 
		s_E108_C1_L				  :std_logic_vector(11 downto 0) := x"0D6"; 
		s_E109_C1_L				  :std_logic_vector(11 downto 0) := x"0D8"; 
		s_E110_C1_L				  :std_logic_vector(11 downto 0) := x"0DA"; 
		s_E111_C1_L				  :std_logic_vector(11 downto 0) := x"0DC"; 
		s_E112_C1_L				  :std_logic_vector(11 downto 0) := x"0DE"; 
		s_E113_C1_L				  :std_logic_vector(11 downto 0) := x"0E0"; 
		s_E114_C1_L				  :std_logic_vector(11 downto 0) := x"0E2"; 
		s_E115_C1_L				  :std_logic_vector(11 downto 0) := x"0E4"; 
		s_E116_C1_L				  :std_logic_vector(11 downto 0) := x"0E6"; 
		s_E117_C1_L				  :std_logic_vector(11 downto 0) := x"0E8"; 
		s_E118_C1_L				  :std_logic_vector(11 downto 0) := x"0EA"; 
		s_E119_C1_L				  :std_logic_vector(11 downto 0) := x"0EC"; 
		s_E120_C1_L				  :std_logic_vector(11 downto 0) := x"0EE"; 
		s_E121_C1_L				  :std_logic_vector(11 downto 0) := x"0F0"; 
		s_E122_C1_L				  :std_logic_vector(11 downto 0) := x"0F2"; 
		s_E123_C1_L				  :std_logic_vector(11 downto 0) := x"0F4"; 
		s_E124_C1_L				  :std_logic_vector(11 downto 0) := x"0F6"; 
		s_E125_C1_L				  :std_logic_vector(11 downto 0) := x"0F8"; 
		s_E126_C1_L				  :std_logic_vector(11 downto 0) := x"0FA"; 
		s_E127_C1_L				  :std_logic_vector(11 downto 0) := x"0FC"; 
		s_E128_C1_L				  :std_logic_vector(11 downto 0) := x"0FE"; 
		s_E129_C1_L				  :std_logic_vector(11 downto 0) := x"100"; 
		s_E130_C1_L				  :std_logic_vector(11 downto 0) := x"102"; 
		s_E131_C1_L				  :std_logic_vector(11 downto 0) := x"104"; 
		s_E132_C1_L				  :std_logic_vector(11 downto 0) := x"106"; 
		s_E133_C1_L				  :std_logic_vector(11 downto 0) := x"108"; 
		s_E134_C1_L				  :std_logic_vector(11 downto 0) := x"10A"; 
		s_E135_C1_L				  :std_logic_vector(11 downto 0) := x"10C"; 
		s_E136_C1_L				  :std_logic_vector(11 downto 0) := x"10E"; 
		s_E137_C1_L				  :std_logic_vector(11 downto 0) := x"110"; 
		s_E138_C1_L				  :std_logic_vector(11 downto 0) := x"112"; 
		s_E139_C1_L				  :std_logic_vector(11 downto 0) := x"114"; 
		s_E140_C1_L				  :std_logic_vector(11 downto 0) := x"116"; 
		s_E141_C1_L				  :std_logic_vector(11 downto 0) := x"118"; 
		s_E142_C1_L				  :std_logic_vector(11 downto 0) := x"11A"; 
		s_E143_C1_L				  :std_logic_vector(11 downto 0) := x"11C"; 
		s_E144_C1_L				  :std_logic_vector(11 downto 0) := x"11E"; 
		s_E145_C1_L				  :std_logic_vector(11 downto 0) := x"120"; 
		s_E146_C1_L				  :std_logic_vector(11 downto 0) := x"122"; 
		s_E147_C1_L				  :std_logic_vector(11 downto 0) := x"124"; 
		s_E148_C1_L				  :std_logic_vector(11 downto 0) := x"126"; 
		s_E149_C1_L				  :std_logic_vector(11 downto 0) := x"128"; 
		s_E150_C1_L				  :std_logic_vector(11 downto 0) := x"12A"; 
		s_E151_C1_L				  :std_logic_vector(11 downto 0) := x"12C"; 
		s_E152_C1_L				  :std_logic_vector(11 downto 0) := x"12E"; 
		s_E153_C1_L				  :std_logic_vector(11 downto 0) := x"130"; 
		s_E154_C1_L				  :std_logic_vector(11 downto 0) := x"132"; 
		s_E155_C1_L				  :std_logic_vector(11 downto 0) := x"134"; 
		s_E156_C1_L				  :std_logic_vector(11 downto 0) := x"136"; 
		s_E157_C1_L				  :std_logic_vector(11 downto 0) := x"138"; 
		s_E158_C1_L				  :std_logic_vector(11 downto 0) := x"13A"; 
		s_E159_C1_L				  :std_logic_vector(11 downto 0) := x"13C"; 
		s_E160_C1_L				  :std_logic_vector(11 downto 0) := x"13E"; 
		s_E161_C1_L				  :std_logic_vector(11 downto 0) := x"140"; 
		s_E162_C1_L				  :std_logic_vector(11 downto 0) := x"142"; 
		s_E163_C1_L				  :std_logic_vector(11 downto 0) := x"144"; 
		s_E164_C1_L				  :std_logic_vector(11 downto 0) := x"146"; 
		s_E165_C1_L				  :std_logic_vector(11 downto 0) := x"148"; 
		s_E166_C1_L				  :std_logic_vector(11 downto 0) := x"14A"; 
		s_E167_C1_L				  :std_logic_vector(11 downto 0) := x"14C"; 
		s_E168_C1_L				  :std_logic_vector(11 downto 0) := x"14E"; 
		s_E169_C1_L				  :std_logic_vector(11 downto 0) := x"150"; 
		s_E170_C1_L				  :std_logic_vector(11 downto 0) := x"152"; 
		s_E171_C1_L				  :std_logic_vector(11 downto 0) := x"154"; 
		s_E172_C1_L				  :std_logic_vector(11 downto 0) := x"156"; 
		s_E173_C1_L				  :std_logic_vector(11 downto 0) := x"158"; 
		s_E174_C1_L				  :std_logic_vector(11 downto 0) := x"15A"; 
		s_E175_C1_L				  :std_logic_vector(11 downto 0) := x"15C"; 
		s_E176_C1_L				  :std_logic_vector(11 downto 0) := x"15E"; 
		s_E177_C1_L				  :std_logic_vector(11 downto 0) := x"160"; 
		s_E178_C1_L				  :std_logic_vector(11 downto 0) := x"162"; 
		s_E179_C1_L				  :std_logic_vector(11 downto 0) := x"164"; 
		s_E180_C1_L				  :std_logic_vector(11 downto 0) := x"166"; 
		s_E181_C1_L				  :std_logic_vector(11 downto 0) := x"168"; 
		s_E182_C1_L				  :std_logic_vector(11 downto 0) := x"16A"; 
		s_E183_C1_L				  :std_logic_vector(11 downto 0) := x"16C"; 
		s_E184_C1_L				  :std_logic_vector(11 downto 0) := x"16E"; 
		s_E185_C1_L				  :std_logic_vector(11 downto 0) := x"170"; 
		s_E186_C1_L				  :std_logic_vector(11 downto 0) := x"172"; 
		s_E187_C1_L				  :std_logic_vector(11 downto 0) := x"174"; 
		s_E188_C1_L				  :std_logic_vector(11 downto 0) := x"176"; 
		s_E189_C1_L				  :std_logic_vector(11 downto 0) := x"178"; 
		s_E190_C1_L				  :std_logic_vector(11 downto 0) := x"17A"; 
		s_E191_C1_L				  :std_logic_vector(11 downto 0) := x"17C"; 
		s_E192_C1_L				  :std_logic_vector(11 downto 0) := x"17E"; 
		s_E193_C1_L				  :std_logic_vector(11 downto 0) := x"180"; 
		s_E194_C1_L				  :std_logic_vector(11 downto 0) := x"182"; 
		s_E195_C1_L				  :std_logic_vector(11 downto 0) := x"184"; 
		s_E196_C1_L				  :std_logic_vector(11 downto 0) := x"186"; 
		s_E197_C1_L				  :std_logic_vector(11 downto 0) := x"188"; 
		s_E198_C1_L				  :std_logic_vector(11 downto 0) := x"18A"; 
		s_E199_C1_L				  :std_logic_vector(11 downto 0) := x"18C"; 
		s_E200_C1_L				  :std_logic_vector(11 downto 0) := x"18E"; 
		s_E201_C1_L				  :std_logic_vector(11 downto 0) := x"190"; 
		s_E202_C1_L				  :std_logic_vector(11 downto 0) := x"192"; 
		s_E203_C1_L				  :std_logic_vector(11 downto 0) := x"194"; 
		s_E204_C1_L				  :std_logic_vector(11 downto 0) := x"196"; 
		s_E205_C1_L				  :std_logic_vector(11 downto 0) := x"198"; 
		s_E206_C1_L				  :std_logic_vector(11 downto 0) := x"19A"; 
		s_E207_C1_L				  :std_logic_vector(11 downto 0) := x"19C"; 
		s_E208_C1_L				  :std_logic_vector(11 downto 0) := x"19E"; 
		s_E209_C1_L				  :std_logic_vector(11 downto 0) := x"1A0"; 
		s_E210_C1_L				  :std_logic_vector(11 downto 0) := x"1A2"; 
		s_E211_C1_L				  :std_logic_vector(11 downto 0) := x"1A4"; 
		s_E212_C1_L				  :std_logic_vector(11 downto 0) := x"1A6"; 
		s_E213_C1_L				  :std_logic_vector(11 downto 0) := x"1A8"; 
		s_E214_C1_L				  :std_logic_vector(11 downto 0) := x"1AA"; 
		s_E215_C1_L				  :std_logic_vector(11 downto 0) := x"1AC"; 
		s_E216_C1_L				  :std_logic_vector(11 downto 0) := x"1AE"; 
		s_E217_C1_L				  :std_logic_vector(11 downto 0) := x"1B0"; 
		s_E218_C1_L				  :std_logic_vector(11 downto 0) := x"1B2"; 
		s_E219_C1_L				  :std_logic_vector(11 downto 0) := x"1B4"; 
		s_E220_C1_L				  :std_logic_vector(11 downto 0) := x"1B6"; 
		s_E221_C1_L				  :std_logic_vector(11 downto 0) := x"1B8"; 
		s_E222_C1_L				  :std_logic_vector(11 downto 0) := x"1BA"; 
		s_E223_C1_L				  :std_logic_vector(11 downto 0) := x"1BC"; 
		s_E224_C1_L				  :std_logic_vector(11 downto 0) := x"1BE"; 
		s_E225_C1_L				  :std_logic_vector(11 downto 0) := x"1C0"; 
		s_E226_C1_L				  :std_logic_vector(11 downto 0) := x"1C2"; 
		s_E227_C1_L				  :std_logic_vector(11 downto 0) := x"1C4"; 
		s_E228_C1_L				  :std_logic_vector(11 downto 0) := x"1C6"; 
		s_E229_C1_L				  :std_logic_vector(11 downto 0) := x"1C8"; 
		s_E230_C1_L				  :std_logic_vector(11 downto 0) := x"1CA"; 
		s_E231_C1_L				  :std_logic_vector(11 downto 0) := x"1CC"; 
		s_E232_C1_L				  :std_logic_vector(11 downto 0) := x"1CE"; 
		s_E233_C1_L				  :std_logic_vector(11 downto 0) := x"1D0"; 
		s_E234_C1_L				  :std_logic_vector(11 downto 0) := x"1D2"; 
		s_E235_C1_L				  :std_logic_vector(11 downto 0) := x"1D4"; 
		s_E236_C1_L				  :std_logic_vector(11 downto 0) := x"1D6"; 
		s_E237_C1_L				  :std_logic_vector(11 downto 0) := x"1D8"; 
		s_E238_C1_L				  :std_logic_vector(11 downto 0) := x"1DA"; 
		s_E239_C1_L				  :std_logic_vector(11 downto 0) := x"1DC"; 
		s_E240_C1_L				  :std_logic_vector(11 downto 0) := x"1DE"; 
		s_E241_C1_L				  :std_logic_vector(11 downto 0) := x"1E0"; 
		s_E242_C1_L				  :std_logic_vector(11 downto 0) := x"1E2"; 
		s_E243_C1_L				  :std_logic_vector(11 downto 0) := x"1E4"; 
		s_E244_C1_L				  :std_logic_vector(11 downto 0) := x"1E6"; 
		s_E245_C1_L				  :std_logic_vector(11 downto 0) := x"1E8"; 
		s_E246_C1_L				  :std_logic_vector(11 downto 0) := x"1EA"; 
		s_E247_C1_L				  :std_logic_vector(11 downto 0) := x"1EC"; 
		s_E248_C1_L				  :std_logic_vector(11 downto 0) := x"1EE"; 
		s_E249_C1_L				  :std_logic_vector(11 downto 0) := x"1F0"; 
		s_E250_C1_L				  :std_logic_vector(11 downto 0) := x"1F2"; 
		s_E251_C1_L				  :std_logic_vector(11 downto 0) := x"1F4"; 
		s_E252_C1_L				  :std_logic_vector(11 downto 0) := x"1F6"; 
		s_E253_C1_L				  :std_logic_vector(11 downto 0) := x"1F8"; 
		s_E254_C1_L				  :std_logic_vector(11 downto 0) := x"1FA"; 
		s_E255_C1_L				  :std_logic_vector(11 downto 0) := x"1FC"; 
		s_E256_C1_L				  :std_logic_vector(11 downto 0) := x"1FE"; 
		s_E257_C1_L				  :std_logic_vector(11 downto 0) := x"200"; 
		s_E258_C1_L				  :std_logic_vector(11 downto 0) := x"202"; 
		s_E259_C1_L				  :std_logic_vector(11 downto 0) := x"204"; 
		s_E260_C1_L				  :std_logic_vector(11 downto 0) := x"206"; 
		s_E261_C1_L				  :std_logic_vector(11 downto 0) := x"208"; 
		s_E262_C1_L				  :std_logic_vector(11 downto 0) := x"20A"; 
		s_E263_C1_L				  :std_logic_vector(11 downto 0) := x"20C"; 
		s_E264_C1_L				  :std_logic_vector(11 downto 0) := x"20E"; 
		s_E265_C1_L				  :std_logic_vector(11 downto 0) := x"210"; 
		s_E266_C1_L				  :std_logic_vector(11 downto 0) := x"212"; 
		s_E267_C1_L				  :std_logic_vector(11 downto 0) := x"214"; 
		s_E268_C1_L				  :std_logic_vector(11 downto 0) := x"216"; 
		s_E269_C1_L				  :std_logic_vector(11 downto 0) := x"218"; 
		s_E270_C1_L				  :std_logic_vector(11 downto 0) := x"21A"; 
		s_E271_C1_L				  :std_logic_vector(11 downto 0) := x"21C"; 
		s_E272_C1_L				  :std_logic_vector(11 downto 0) := x"21E"; 
		s_E273_C1_L				  :std_logic_vector(11 downto 0) := x"220"; 
		s_E274_C1_L				  :std_logic_vector(11 downto 0) := x"222"; 
		s_E275_C1_L				  :std_logic_vector(11 downto 0) := x"224"; 
		s_E276_C1_L				  :std_logic_vector(11 downto 0) := x"226"; 
		s_E277_C1_L				  :std_logic_vector(11 downto 0) := x"228"; 
		s_E278_C1_L				  :std_logic_vector(11 downto 0) := x"22A"; 
		s_E279_C1_L				  :std_logic_vector(11 downto 0) := x"22C"; 
		s_E280_C1_L				  :std_logic_vector(11 downto 0) := x"22E"; 
		s_E281_C1_L				  :std_logic_vector(11 downto 0) := x"230"; 
		s_E282_C1_L				  :std_logic_vector(11 downto 0) := x"232"; 
		s_E283_C1_L				  :std_logic_vector(11 downto 0) := x"234"; 
		s_E284_C1_L				  :std_logic_vector(11 downto 0) := x"236"; 
		s_E285_C1_L				  :std_logic_vector(11 downto 0) := x"238"; 
		s_E286_C1_L				  :std_logic_vector(11 downto 0) := x"23A"; 
		s_E287_C1_L				  :std_logic_vector(11 downto 0) := x"23C"; 
		s_E288_C1_L				  :std_logic_vector(11 downto 0) := x"23E"; 
		s_E289_C1_L				  :std_logic_vector(11 downto 0) := x"240"; 
		s_E290_C1_L				  :std_logic_vector(11 downto 0) := x"242"; 
		s_E291_C1_L				  :std_logic_vector(11 downto 0) := x"244"; 
		s_E292_C1_L				  :std_logic_vector(11 downto 0) := x"246"; 
		s_E293_C1_L				  :std_logic_vector(11 downto 0) := x"248"; 
		s_E294_C1_L				  :std_logic_vector(11 downto 0) := x"24A"; 
		s_E295_C1_L				  :std_logic_vector(11 downto 0) := x"24C"; 
		s_E296_C1_L				  :std_logic_vector(11 downto 0) := x"24E"; 
		s_E297_C1_L				  :std_logic_vector(11 downto 0) := x"250"; 
		s_E298_C1_L				  :std_logic_vector(11 downto 0) := x"252"; 
		s_E299_C1_L				  :std_logic_vector(11 downto 0) := x"254"; 
		s_E300_C1_L				  :std_logic_vector(11 downto 0) := x"256"; 
		s_E301_C1_L				  :std_logic_vector(11 downto 0) := x"258"; 
		s_E302_C1_L				  :std_logic_vector(11 downto 0) := x"25A"; 
		s_E303_C1_L				  :std_logic_vector(11 downto 0) := x"25C"; 
		s_E304_C1_L				  :std_logic_vector(11 downto 0) := x"25E"; 
		s_E305_C1_L				  :std_logic_vector(11 downto 0) := x"260"; 
		s_E306_C1_L				  :std_logic_vector(11 downto 0) := x"262"; 
		s_E307_C1_L				  :std_logic_vector(11 downto 0) := x"264"; 
		s_E308_C1_L				  :std_logic_vector(11 downto 0) := x"266"; 
		s_E309_C1_L				  :std_logic_vector(11 downto 0) := x"268"; 
		s_E310_C1_L				  :std_logic_vector(11 downto 0) := x"26A"; 
		s_E311_C1_L				  :std_logic_vector(11 downto 0) := x"26C"; 
		s_E312_C1_L				  :std_logic_vector(11 downto 0) := x"26E"; 
		s_E313_C1_L				  :std_logic_vector(11 downto 0) := x"270"; 
		s_E314_C1_L				  :std_logic_vector(11 downto 0) := x"272"; 
		s_E315_C1_L				  :std_logic_vector(11 downto 0) := x"274"; 
		s_E316_C1_L				  :std_logic_vector(11 downto 0) := x"276"; 
		s_E317_C1_L				  :std_logic_vector(11 downto 0) := x"278"; 
		s_E318_C1_L				  :std_logic_vector(11 downto 0) := x"27A"; 
		s_E319_C1_L				  :std_logic_vector(11 downto 0) := x"27C"; 
		s_E320_C1_L				  :std_logic_vector(11 downto 0) := x"27E"; 
		s_E321_C1_L				  :std_logic_vector(11 downto 0) := x"280"; 
		s_E322_C1_L				  :std_logic_vector(11 downto 0) := x"282"; 
		s_E323_C1_L				  :std_logic_vector(11 downto 0) := x"284"; 
		s_E324_C1_L				  :std_logic_vector(11 downto 0) := x"286"; 
		s_E325_C1_L				  :std_logic_vector(11 downto 0) := x"288"; 
		s_E326_C1_L				  :std_logic_vector(11 downto 0) := x"28A"; 
		s_E327_C1_L				  :std_logic_vector(11 downto 0) := x"28C"; 
		s_E328_C1_L				  :std_logic_vector(11 downto 0) := x"28E"; 
		s_E329_C1_L				  :std_logic_vector(11 downto 0) := x"290"; 
		s_E330_C1_L				  :std_logic_vector(11 downto 0) := x"292"; 
		s_E331_C1_L				  :std_logic_vector(11 downto 0) := x"294"; 
		s_E332_C1_L				  :std_logic_vector(11 downto 0) := x"296"; 
		s_E333_C1_L				  :std_logic_vector(11 downto 0) := x"298"; 
		s_E334_C1_L				  :std_logic_vector(11 downto 0) := x"29A"; 
		s_E335_C1_L				  :std_logic_vector(11 downto 0) := x"29C"; 
		s_E336_C1_L				  :std_logic_vector(11 downto 0) := x"29E"; 
		s_E337_C1_L				  :std_logic_vector(11 downto 0) := x"2A0"; 
		s_E338_C1_L				  :std_logic_vector(11 downto 0) := x"2A2"; 
		s_E339_C1_L				  :std_logic_vector(11 downto 0) := x"2A4"; 
		s_E340_C1_L				  :std_logic_vector(11 downto 0) := x"2A6"; 
		s_E341_C1_L				  :std_logic_vector(11 downto 0) := x"2A8"; 
		s_E342_C1_L				  :std_logic_vector(11 downto 0) := x"2AA"; 
		s_E343_C1_L				  :std_logic_vector(11 downto 0) := x"2AC"; 
		s_E344_C1_L				  :std_logic_vector(11 downto 0) := x"2AE"; 
		s_E345_C1_L				  :std_logic_vector(11 downto 0) := x"2B0"; 
		s_E346_C1_L				  :std_logic_vector(11 downto 0) := x"2B2"; 
		s_E347_C1_L				  :std_logic_vector(11 downto 0) := x"2B4"; 
		s_E348_C1_L				  :std_logic_vector(11 downto 0) := x"2B6"; 
		s_E349_C1_L				  :std_logic_vector(11 downto 0) := x"2B8"; 
		s_E350_C1_L				  :std_logic_vector(11 downto 0) := x"2BA"; 
		s_E351_C1_L				  :std_logic_vector(11 downto 0) := x"2BC"; 
		s_E352_C1_L				  :std_logic_vector(11 downto 0) := x"2BE"; 
		s_E353_C1_L				  :std_logic_vector(11 downto 0) := x"2C0"; 
		s_E354_C1_L				  :std_logic_vector(11 downto 0) := x"2C2"; 
		s_E355_C1_L				  :std_logic_vector(11 downto 0) := x"2C4"; 
		s_E356_C1_L				  :std_logic_vector(11 downto 0) := x"2C6"; 
		s_E357_C1_L				  :std_logic_vector(11 downto 0) := x"2C8"; 
		s_E358_C1_L				  :std_logic_vector(11 downto 0) := x"2CA"; 
		s_E359_C1_L				  :std_logic_vector(11 downto 0) := x"2CC"; 
		s_E360_C1_L				  :std_logic_vector(11 downto 0) := x"2CE"; 
		s_E361_C1_L				  :std_logic_vector(11 downto 0) := x"2D0"; 
		s_E362_C1_L				  :std_logic_vector(11 downto 0) := x"2D2"; 
		s_E363_C1_L				  :std_logic_vector(11 downto 0) := x"2D4"; 
		s_E364_C1_L				  :std_logic_vector(11 downto 0) := x"2D6"; 
		s_E365_C1_L				  :std_logic_vector(11 downto 0) := x"2D8"; 
		s_E366_C1_L				  :std_logic_vector(11 downto 0) := x"2DA"; 
		s_E367_C1_L				  :std_logic_vector(11 downto 0) := x"2DC"; 
		s_E368_C1_L				  :std_logic_vector(11 downto 0) := x"2DE"; 
		s_E369_C1_L				  :std_logic_vector(11 downto 0) := x"2E0"; 
		s_E370_C1_L				  :std_logic_vector(11 downto 0) := x"2E2"; 
		s_E371_C1_L				  :std_logic_vector(11 downto 0) := x"2E4"; 
		s_E372_C1_L				  :std_logic_vector(11 downto 0) := x"2E6"; 
		s_E373_C1_L				  :std_logic_vector(11 downto 0) := x"2E8"; 
		s_E374_C1_L				  :std_logic_vector(11 downto 0) := x"2EA"; 
		s_E375_C1_L				  :std_logic_vector(11 downto 0) := x"2EC"; 
		s_E376_C1_L				  :std_logic_vector(11 downto 0) := x"2EE"; 
		s_E377_C1_L				  :std_logic_vector(11 downto 0) := x"2F0"; 
		s_E378_C1_L				  :std_logic_vector(11 downto 0) := x"2F2"; 
		s_E379_C1_L				  :std_logic_vector(11 downto 0) := x"2F4"; 
		s_E380_C1_L				  :std_logic_vector(11 downto 0) := x"2F6"; 
		s_E381_C1_L				  :std_logic_vector(11 downto 0) := x"2F8"; 
		s_E382_C1_L				  :std_logic_vector(11 downto 0) := x"2FA"; 
		s_E383_C1_L				  :std_logic_vector(11 downto 0) := x"2FC"; 
		s_E384_C1_L				  :std_logic_vector(11 downto 0) := x"2FE"; 
		s_E385_C1_L				  :std_logic_vector(11 downto 0) := x"300"; 
		s_E386_C1_L				  :std_logic_vector(11 downto 0) := x"302"; 
		s_E387_C1_L				  :std_logic_vector(11 downto 0) := x"304"; 
		s_E388_C1_L				  :std_logic_vector(11 downto 0) := x"306"; 
		s_E389_C1_L				  :std_logic_vector(11 downto 0) := x"308"; 
		s_E390_C1_L				  :std_logic_vector(11 downto 0) := x"30A"; 
		s_E391_C1_L				  :std_logic_vector(11 downto 0) := x"30C"; 
		s_E392_C1_L				  :std_logic_vector(11 downto 0) := x"30E"; 
		s_E393_C1_L				  :std_logic_vector(11 downto 0) := x"310"; 
		s_E394_C1_L				  :std_logic_vector(11 downto 0) := x"312"; 
		s_E395_C1_L				  :std_logic_vector(11 downto 0) := x"314"; 
		s_E396_C1_L				  :std_logic_vector(11 downto 0) := x"316"; 
		s_E397_C1_L				  :std_logic_vector(11 downto 0) := x"318"; 
		s_E398_C1_L				  :std_logic_vector(11 downto 0) := x"31A"; 
		s_E399_C1_L				  :std_logic_vector(11 downto 0) := x"31C"; 
		s_E400_C1_L				  :std_logic_vector(11 downto 0) := x"31E"; 
		s_E401_C1_L				  :std_logic_vector(11 downto 0) := x"320"; 
		s_E402_C1_L				  :std_logic_vector(11 downto 0) := x"322"; 
		s_E403_C1_L				  :std_logic_vector(11 downto 0) := x"324"; 
		s_E404_C1_L				  :std_logic_vector(11 downto 0) := x"326"; 
		s_E405_C1_L				  :std_logic_vector(11 downto 0) := x"328"; 
		s_E406_C1_L				  :std_logic_vector(11 downto 0) := x"32A"; 
		s_E407_C1_L				  :std_logic_vector(11 downto 0) := x"32C"; 
		s_E408_C1_L				  :std_logic_vector(11 downto 0) := x"32E"; 
		s_E409_C1_L				  :std_logic_vector(11 downto 0) := x"330"; 
		s_E410_C1_L				  :std_logic_vector(11 downto 0) := x"332"; 
		s_E411_C1_L				  :std_logic_vector(11 downto 0) := x"334"; 
		s_E412_C1_L				  :std_logic_vector(11 downto 0) := x"336"; 
		s_E413_C1_L				  :std_logic_vector(11 downto 0) := x"338"; 
		s_E414_C1_L				  :std_logic_vector(11 downto 0) := x"33A"; 
		s_E415_C1_L				  :std_logic_vector(11 downto 0) := x"33C"; 
		s_E416_C1_L				  :std_logic_vector(11 downto 0) := x"33E"; 
		s_E417_C1_L				  :std_logic_vector(11 downto 0) := x"340"; 
		s_E418_C1_L				  :std_logic_vector(11 downto 0) := x"342"; 
		s_E419_C1_L				  :std_logic_vector(11 downto 0) := x"344"; 
		s_E420_C1_L				  :std_logic_vector(11 downto 0) := x"346"; 
		s_E421_C1_L				  :std_logic_vector(11 downto 0) := x"348"; 
		s_E422_C1_L				  :std_logic_vector(11 downto 0) := x"34A"; 
		s_E423_C1_L				  :std_logic_vector(11 downto 0) := x"34C"; 
		s_E424_C1_L				  :std_logic_vector(11 downto 0) := x"34E"; 
		s_E425_C1_L				  :std_logic_vector(11 downto 0) := x"350"; 
		s_E426_C1_L				  :std_logic_vector(11 downto 0) := x"352"; 
		s_E427_C1_L				  :std_logic_vector(11 downto 0) := x"354"; 
		s_E428_C1_L				  :std_logic_vector(11 downto 0) := x"356"; 
		s_E429_C1_L				  :std_logic_vector(11 downto 0) := x"358"; 
		s_E430_C1_L				  :std_logic_vector(11 downto 0) := x"35A"; 
		s_E431_C1_L				  :std_logic_vector(11 downto 0) := x"35C"; 
		s_E432_C1_L				  :std_logic_vector(11 downto 0) := x"35E"; 
		s_E433_C1_L				  :std_logic_vector(11 downto 0) := x"360"; 
		s_E434_C1_L				  :std_logic_vector(11 downto 0) := x"362"; 
		s_E435_C1_L				  :std_logic_vector(11 downto 0) := x"364"; 
		s_E436_C1_L				  :std_logic_vector(11 downto 0) := x"366"; 
		s_E437_C1_L				  :std_logic_vector(11 downto 0) := x"368"; 
		s_E438_C1_L				  :std_logic_vector(11 downto 0) := x"36A"; 
		s_E439_C1_L				  :std_logic_vector(11 downto 0) := x"36C"; 
		s_E440_C1_L				  :std_logic_vector(11 downto 0) := x"36E"; 
		s_E441_C1_L				  :std_logic_vector(11 downto 0) := x"370"; 
		s_E442_C1_L				  :std_logic_vector(11 downto 0) := x"372"; 
		s_E443_C1_L				  :std_logic_vector(11 downto 0) := x"374"; 
		s_E444_C1_L				  :std_logic_vector(11 downto 0) := x"376"; 
		s_E445_C1_L				  :std_logic_vector(11 downto 0) := x"378"; 
		s_E446_C1_L				  :std_logic_vector(11 downto 0) := x"37A"; 
		s_E447_C1_L				  :std_logic_vector(11 downto 0) := x"37C"; 
		s_E448_C1_L				  :std_logic_vector(11 downto 0) := x"37E"; 
		s_E449_C1_L				  :std_logic_vector(11 downto 0) := x"380"; 
		s_E450_C1_L				  :std_logic_vector(11 downto 0) := x"382"; 
		s_E451_C1_L				  :std_logic_vector(11 downto 0) := x"384"; 
		s_E452_C1_L				  :std_logic_vector(11 downto 0) := x"386"; 
		s_E453_C1_L				  :std_logic_vector(11 downto 0) := x"388"; 
		s_E454_C1_L				  :std_logic_vector(11 downto 0) := x"38A"; 
		s_E455_C1_L				  :std_logic_vector(11 downto 0) := x"38C"; 
		s_E456_C1_L				  :std_logic_vector(11 downto 0) := x"38E"; 
		s_E457_C1_L				  :std_logic_vector(11 downto 0) := x"390"; 
		s_E458_C1_L				  :std_logic_vector(11 downto 0) := x"392"; 
		s_E459_C1_L				  :std_logic_vector(11 downto 0) := x"394"; 
		s_E460_C1_L				  :std_logic_vector(11 downto 0) := x"396"; 
		s_E461_C1_L				  :std_logic_vector(11 downto 0) := x"398"; 
		s_E462_C1_L				  :std_logic_vector(11 downto 0) := x"39A"; 
		s_E463_C1_L				  :std_logic_vector(11 downto 0) := x"39C"; 
		s_E464_C1_L				  :std_logic_vector(11 downto 0) := x"39E"; 
		s_E465_C1_L				  :std_logic_vector(11 downto 0) := x"3A0"; 
		s_E466_C1_L				  :std_logic_vector(11 downto 0) := x"3A2"; 
		s_E467_C1_L				  :std_logic_vector(11 downto 0) := x"3A4"; 
		s_E468_C1_L				  :std_logic_vector(11 downto 0) := x"3A6"; 
		s_E469_C1_L				  :std_logic_vector(11 downto 0) := x"3A8"; 
		s_E470_C1_L				  :std_logic_vector(11 downto 0) := x"3AA"; 
		s_E471_C1_L				  :std_logic_vector(11 downto 0) := x"3AC"; 
		s_E472_C1_L				  :std_logic_vector(11 downto 0) := x"3AE"; 
		s_E473_C1_L				  :std_logic_vector(11 downto 0) := x"3B0"; 
		s_E474_C1_L				  :std_logic_vector(11 downto 0) := x"3B2"; 
		s_E475_C1_L				  :std_logic_vector(11 downto 0) := x"3B4"; 
		s_E476_C1_L				  :std_logic_vector(11 downto 0) := x"3B6"; 
		s_E477_C1_L				  :std_logic_vector(11 downto 0) := x"3B8"; 
		s_E478_C1_L				  :std_logic_vector(11 downto 0) := x"3BA"; 
		s_E479_C1_L				  :std_logic_vector(11 downto 0) := x"3BC"; 
		s_E480_C1_L				  :std_logic_vector(11 downto 0) := x"3BE"; 
		s_E481_C1_L				  :std_logic_vector(11 downto 0) := x"3C0"; 
		s_E482_C1_L				  :std_logic_vector(11 downto 0) := x"3C2"; 
		s_E483_C1_L				  :std_logic_vector(11 downto 0) := x"3C4"; 
		s_E484_C1_L				  :std_logic_vector(11 downto 0) := x"3C6"; 
		s_E485_C1_L				  :std_logic_vector(11 downto 0) := x"3C8"; 
		s_E486_C1_L				  :std_logic_vector(11 downto 0) := x"3CA"; 
		s_E487_C1_L				  :std_logic_vector(11 downto 0) := x"3CC"; 
		s_E488_C1_L				  :std_logic_vector(11 downto 0) := x"3CE"; 
		s_E489_C1_L				  :std_logic_vector(11 downto 0) := x"3D0"; 
		s_E490_C1_L				  :std_logic_vector(11 downto 0) := x"3D2"; 
		s_E491_C1_L				  :std_logic_vector(11 downto 0) := x"3D4"; 
		s_E492_C1_L				  :std_logic_vector(11 downto 0) := x"3D6"; 
		s_E493_C1_L				  :std_logic_vector(11 downto 0) := x"3D8"; 
		s_E494_C1_L				  :std_logic_vector(11 downto 0) := x"3DA"; 
		s_E495_C1_L				  :std_logic_vector(11 downto 0) := x"3DC"; 
		s_E496_C1_L				  :std_logic_vector(11 downto 0) := x"3DE"; 
		s_E497_C1_L				  :std_logic_vector(11 downto 0) := x"3E0"; 
		s_E498_C1_L				  :std_logic_vector(11 downto 0) := x"3E2"; 
		s_E499_C1_L				  :std_logic_vector(11 downto 0) := x"3E4"; 
		s_E500_C1_L				  :std_logic_vector(11 downto 0) := x"3E6"; 
		s_E501_C1_L				  :std_logic_vector(11 downto 0) := x"3E8"; 
		s_E502_C1_L				  :std_logic_vector(11 downto 0) := x"3EA"; 
		s_E503_C1_L				  :std_logic_vector(11 downto 0) := x"3EC"; 
		s_E504_C1_L				  :std_logic_vector(11 downto 0) := x"3EE"; 
		s_E505_C1_L				  :std_logic_vector(11 downto 0) := x"3F0"; 
		s_E506_C1_L				  :std_logic_vector(11 downto 0) := x"3F2"; 
		s_E507_C1_L				  :std_logic_vector(11 downto 0) := x"3F4"; 
		s_E508_C1_L				  :std_logic_vector(11 downto 0) := x"3F6"; 
		s_E509_C1_L				  :std_logic_vector(11 downto 0) := x"3F8"; 
		s_E510_C1_L				  :std_logic_vector(11 downto 0) := x"3FA"; 
		s_E511_C1_L				  :std_logic_vector(11 downto 0) := x"3FC"; 
		s_E512_C1_L				  :std_logic_vector(11 downto 0) := x"3FE"; 
		s_E513_C1_L				  :std_logic_vector(11 downto 0) := x"400"; 
		s_E514_C1_L				  :std_logic_vector(11 downto 0) := x"402"; 
		s_E515_C1_L				  :std_logic_vector(11 downto 0) := x"404"; 
		s_E516_C1_L				  :std_logic_vector(11 downto 0) := x"406"; 
		s_E517_C1_L				  :std_logic_vector(11 downto 0) := x"408"; 
		s_E518_C1_L				  :std_logic_vector(11 downto 0) := x"40A"; 
		s_E519_C1_L				  :std_logic_vector(11 downto 0) := x"40C"; 
		s_E520_C1_L				  :std_logic_vector(11 downto 0) := x"40E"; 
		s_E521_C1_L				  :std_logic_vector(11 downto 0) := x"410"; 
		s_E522_C1_L				  :std_logic_vector(11 downto 0) := x"412"; 
		s_E523_C1_L				  :std_logic_vector(11 downto 0) := x"414"; 
		s_E524_C1_L				  :std_logic_vector(11 downto 0) := x"416"; 
		s_E525_C1_L				  :std_logic_vector(11 downto 0) := x"418"; 
		s_E526_C1_L				  :std_logic_vector(11 downto 0) := x"41A"; 
		s_E527_C1_L				  :std_logic_vector(11 downto 0) := x"41C"; 
		s_E528_C1_L				  :std_logic_vector(11 downto 0) := x"41E"; 
		s_E529_C1_L				  :std_logic_vector(11 downto 0) := x"420"; 
		s_E530_C1_L				  :std_logic_vector(11 downto 0) := x"422"; 
		s_E531_C1_L				  :std_logic_vector(11 downto 0) := x"424"; 
		s_E532_C1_L				  :std_logic_vector(11 downto 0) := x"426"; 
		s_E533_C1_L				  :std_logic_vector(11 downto 0) := x"428"; 
		s_E534_C1_L				  :std_logic_vector(11 downto 0) := x"42A"; 
		s_E535_C1_L				  :std_logic_vector(11 downto 0) := x"42C"; 
		s_E536_C1_L				  :std_logic_vector(11 downto 0) := x"42E"; 
		s_E537_C1_L				  :std_logic_vector(11 downto 0) := x"430"; 
		s_E538_C1_L				  :std_logic_vector(11 downto 0) := x"432"; 
		s_E539_C1_L				  :std_logic_vector(11 downto 0) := x"434"; 
		s_E540_C1_L				  :std_logic_vector(11 downto 0) := x"436"; 
		s_E541_C1_L				  :std_logic_vector(11 downto 0) := x"438"; 
		s_E542_C1_L				  :std_logic_vector(11 downto 0) := x"43A"; 
		s_E543_C1_L				  :std_logic_vector(11 downto 0) := x"43C"; 
		s_E544_C1_L				  :std_logic_vector(11 downto 0) := x"43E"; 
		s_E545_C1_L				  :std_logic_vector(11 downto 0) := x"440"; 
		s_E546_C1_L				  :std_logic_vector(11 downto 0) := x"442"; 
		s_E547_C1_L				  :std_logic_vector(11 downto 0) := x"444"; 
		s_E548_C1_L				  :std_logic_vector(11 downto 0) := x"446"; 
		s_E549_C1_L				  :std_logic_vector(11 downto 0) := x"448"; 
		s_E550_C1_L				  :std_logic_vector(11 downto 0) := x"44A"; 
		s_E551_C1_L				  :std_logic_vector(11 downto 0) := x"44C"; 
		s_E552_C1_L				  :std_logic_vector(11 downto 0) := x"44E"; 
		s_E553_C1_L				  :std_logic_vector(11 downto 0) := x"450"; 
		s_E554_C1_L				  :std_logic_vector(11 downto 0) := x"452"; 
		s_E555_C1_L				  :std_logic_vector(11 downto 0) := x"454"; 
		s_E556_C1_L				  :std_logic_vector(11 downto 0) := x"456"; 
		s_E557_C1_L				  :std_logic_vector(11 downto 0) := x"458"; 
		s_E558_C1_L				  :std_logic_vector(11 downto 0) := x"45A"; 
		s_E559_C1_L				  :std_logic_vector(11 downto 0) := x"45C"; 
		s_E560_C1_L				  :std_logic_vector(11 downto 0) := x"45E"; 
		s_E561_C1_L				  :std_logic_vector(11 downto 0) := x"460"; 
		s_E562_C1_L				  :std_logic_vector(11 downto 0) := x"462"; 
		s_E563_C1_L				  :std_logic_vector(11 downto 0) := x"464"; 
		s_E564_C1_L				  :std_logic_vector(11 downto 0) := x"466"; 
		s_E565_C1_L				  :std_logic_vector(11 downto 0) := x"468"; 
		s_E566_C1_L				  :std_logic_vector(11 downto 0) := x"46A"; 
		s_E567_C1_L				  :std_logic_vector(11 downto 0) := x"46C"; 
		s_E568_C1_L				  :std_logic_vector(11 downto 0) := x"46E"; 
		s_E569_C1_L				  :std_logic_vector(11 downto 0) := x"470"; 
		s_E570_C1_L				  :std_logic_vector(11 downto 0) := x"472"; 
		s_E571_C1_L				  :std_logic_vector(11 downto 0) := x"474"; 
		s_E572_C1_L				  :std_logic_vector(11 downto 0) := x"476"; 
		s_E573_C1_L				  :std_logic_vector(11 downto 0) := x"478"; 
		s_E574_C1_L				  :std_logic_vector(11 downto 0) := x"47A"; 
		s_E575_C1_L				  :std_logic_vector(11 downto 0) := x"47C"; 
		s_E576_C1_L				  :std_logic_vector(11 downto 0) := x"47E"; 
		s_E577_C1_L				  :std_logic_vector(11 downto 0) := x"480"; 
		s_E578_C1_L				  :std_logic_vector(11 downto 0) := x"482"; 
		s_E579_C1_L				  :std_logic_vector(11 downto 0) := x"484"; 
		s_E580_C1_L				  :std_logic_vector(11 downto 0) := x"486"; 
		s_E581_C1_L				  :std_logic_vector(11 downto 0) := x"488"; 
		s_E582_C1_L				  :std_logic_vector(11 downto 0) := x"48A"; 
		s_E583_C1_L				  :std_logic_vector(11 downto 0) := x"48C"; 
		s_E584_C1_L				  :std_logic_vector(11 downto 0) := x"48E"; 
		s_E585_C1_L				  :std_logic_vector(11 downto 0) := x"490"; 
		s_E586_C1_L				  :std_logic_vector(11 downto 0) := x"492"; 
		s_E587_C1_L				  :std_logic_vector(11 downto 0) := x"494"; 
		s_E588_C1_L				  :std_logic_vector(11 downto 0) := x"496"; 
		s_E589_C1_L				  :std_logic_vector(11 downto 0) := x"498"; 
		s_E590_C1_L				  :std_logic_vector(11 downto 0) := x"49A"; 
		s_E591_C1_L				  :std_logic_vector(11 downto 0) := x"49C"; 
		s_E592_C1_L				  :std_logic_vector(11 downto 0) := x"49E"; 
		s_E593_C1_L				  :std_logic_vector(11 downto 0) := x"4A0"; 
		s_E594_C1_L				  :std_logic_vector(11 downto 0) := x"4A2"; 
		s_E595_C1_L				  :std_logic_vector(11 downto 0) := x"4A4"; 
		s_E596_C1_L				  :std_logic_vector(11 downto 0) := x"4A6"; 
		s_E597_C1_L				  :std_logic_vector(11 downto 0) := x"4A8"; 
		s_E598_C1_L				  :std_logic_vector(11 downto 0) := x"4AA"; 
		s_E599_C1_L				  :std_logic_vector(11 downto 0) := x"4AC"; 
		s_E600_C1_L				  :std_logic_vector(11 downto 0) := x"4AE"; 
		s_E601_C1_L				  :std_logic_vector(11 downto 0) := x"4B0"; 
		s_E602_C1_L				  :std_logic_vector(11 downto 0) := x"4B2"; 
		s_E603_C1_L				  :std_logic_vector(11 downto 0) := x"4B4"; 
		s_E604_C1_L				  :std_logic_vector(11 downto 0) := x"4B6"; 
		s_E605_C1_L				  :std_logic_vector(11 downto 0) := x"4B8"; 
		s_E606_C1_L				  :std_logic_vector(11 downto 0) := x"4BA"; 
		s_E607_C1_L				  :std_logic_vector(11 downto 0) := x"4BC"; 
		s_E608_C1_L				  :std_logic_vector(11 downto 0) := x"4BE"; 
		s_E609_C1_L				  :std_logic_vector(11 downto 0) := x"4C0"; 
		s_E610_C1_L				  :std_logic_vector(11 downto 0) := x"4C2"; 
		s_E611_C1_L				  :std_logic_vector(11 downto 0) := x"4C4"; 
		s_E612_C1_L				  :std_logic_vector(11 downto 0) := x"4C6"; 
		s_E613_C1_L				  :std_logic_vector(11 downto 0) := x"4C8"; 
		s_E614_C1_L				  :std_logic_vector(11 downto 0) := x"4CA"; 
		s_E615_C1_L				  :std_logic_vector(11 downto 0) := x"4CC"; 
		s_E616_C1_L				  :std_logic_vector(11 downto 0) := x"4CE"; 
		s_E617_C1_L				  :std_logic_vector(11 downto 0) := x"4D0"; 
		s_E618_C1_L				  :std_logic_vector(11 downto 0) := x"4D2"; 
		s_E619_C1_L				  :std_logic_vector(11 downto 0) := x"4D4"; 
		s_E620_C1_L				  :std_logic_vector(11 downto 0) := x"4D6"; 
		s_E621_C1_L				  :std_logic_vector(11 downto 0) := x"4D8"; 
		s_E622_C1_L				  :std_logic_vector(11 downto 0) := x"4DA"; 
		s_E623_C1_L				  :std_logic_vector(11 downto 0) := x"4DC"; 
		s_E624_C1_L				  :std_logic_vector(11 downto 0) := x"4DE"; 
		s_E625_C1_L				  :std_logic_vector(11 downto 0) := x"4E0"; 
		s_E626_C1_L				  :std_logic_vector(11 downto 0) := x"4E2"; 
		s_E627_C1_L				  :std_logic_vector(11 downto 0) := x"4E4"; 
		s_E628_C1_L				  :std_logic_vector(11 downto 0) := x"4E6"; 
		s_E629_C1_L				  :std_logic_vector(11 downto 0) := x"4E8"; 
		s_E630_C1_L				  :std_logic_vector(11 downto 0) := x"4EA"; 
		s_E631_C1_L				  :std_logic_vector(11 downto 0) := x"4EC"; 
		s_E632_C1_L				  :std_logic_vector(11 downto 0) := x"4EE"; 
		s_E633_C1_L				  :std_logic_vector(11 downto 0) := x"4F0"; 
		s_E634_C1_L				  :std_logic_vector(11 downto 0) := x"4F2"; 
		s_E635_C1_L				  :std_logic_vector(11 downto 0) := x"4F4"; 
		s_E636_C1_L				  :std_logic_vector(11 downto 0) := x"4F6"; 
		s_E637_C1_L				  :std_logic_vector(11 downto 0) := x"4F8"; 
		s_E638_C1_L				  :std_logic_vector(11 downto 0) := x"4FA"; 
		s_E639_C1_L				  :std_logic_vector(11 downto 0) := x"4FC"; 
		s_E640_C1_L				  :std_logic_vector(11 downto 0) := x"4FE"; 
		s_E641_C1_L				  :std_logic_vector(11 downto 0) := x"500"; 
		s_E642_C1_L				  :std_logic_vector(11 downto 0) := x"502"; 
		s_E643_C1_L				  :std_logic_vector(11 downto 0) := x"504"; 
		s_E644_C1_L				  :std_logic_vector(11 downto 0) := x"506"; 
		s_E645_C1_L				  :std_logic_vector(11 downto 0) := x"508"; 
		s_E646_C1_L				  :std_logic_vector(11 downto 0) := x"50A"; 
		s_E647_C1_L				  :std_logic_vector(11 downto 0) := x"50C"; 
		s_E648_C1_L				  :std_logic_vector(11 downto 0) := x"50E"; 
		s_E649_C1_L				  :std_logic_vector(11 downto 0) := x"510"; 
		s_E650_C1_L				  :std_logic_vector(11 downto 0) := x"512"; 
		s_E651_C1_L				  :std_logic_vector(11 downto 0) := x"514"; 
		s_E652_C1_L				  :std_logic_vector(11 downto 0) := x"516"; 
		s_E653_C1_L				  :std_logic_vector(11 downto 0) := x"518"; 
		s_E654_C1_L				  :std_logic_vector(11 downto 0) := x"51A"; 
		s_E655_C1_L				  :std_logic_vector(11 downto 0) := x"51C"; 
		s_E656_C1_L				  :std_logic_vector(11 downto 0) := x"51E"; 
		s_E657_C1_L				  :std_logic_vector(11 downto 0) := x"520"; 
		s_E658_C1_L				  :std_logic_vector(11 downto 0) := x"522"; 
		s_E659_C1_L				  :std_logic_vector(11 downto 0) := x"524"; 
		s_E660_C1_L				  :std_logic_vector(11 downto 0) := x"526"; 
		s_E661_C1_L				  :std_logic_vector(11 downto 0) := x"528"; 
		s_E662_C1_L				  :std_logic_vector(11 downto 0) := x"52A"; 
		s_E663_C1_L				  :std_logic_vector(11 downto 0) := x"52C"; 
		s_E664_C1_L				  :std_logic_vector(11 downto 0) := x"52E"; 
		s_E665_C1_L				  :std_logic_vector(11 downto 0) := x"530"; 
		s_E666_C1_L				  :std_logic_vector(11 downto 0) := x"532"; 
		s_E667_C1_L				  :std_logic_vector(11 downto 0) := x"534"; 
		s_E668_C1_L				  :std_logic_vector(11 downto 0) := x"536"; 
		s_E669_C1_L				  :std_logic_vector(11 downto 0) := x"538"; 
		s_E670_C1_L				  :std_logic_vector(11 downto 0) := x"53A"; 
		s_E671_C1_L				  :std_logic_vector(11 downto 0) := x"53C"; 
		s_E672_C1_L				  :std_logic_vector(11 downto 0) := x"53E"; 
		s_E673_C1_L				  :std_logic_vector(11 downto 0) := x"540"; 
		s_E674_C1_L				  :std_logic_vector(11 downto 0) := x"542"; 
		s_E675_C1_L				  :std_logic_vector(11 downto 0) := x"544"; 
		s_E676_C1_L				  :std_logic_vector(11 downto 0) := x"546"; 
		s_E677_C1_L				  :std_logic_vector(11 downto 0) := x"548"; 
		s_E678_C1_L				  :std_logic_vector(11 downto 0) := x"54A"; 
		s_E679_C1_L				  :std_logic_vector(11 downto 0) := x"54C"; 
		s_E680_C1_L				  :std_logic_vector(11 downto 0) := x"54E"; 
		s_E681_C1_L				  :std_logic_vector(11 downto 0) := x"550"; 
		s_E682_C1_L				  :std_logic_vector(11 downto 0) := x"552"; 
		s_E683_C1_L				  :std_logic_vector(11 downto 0) := x"554"; 
		s_E684_C1_L				  :std_logic_vector(11 downto 0) := x"556"; 
		s_E685_C1_L				  :std_logic_vector(11 downto 0) := x"558"; 
		s_E686_C1_L				  :std_logic_vector(11 downto 0) := x"55A"; 
		s_E687_C1_L				  :std_logic_vector(11 downto 0) := x"55C"; 
		s_E688_C1_L				  :std_logic_vector(11 downto 0) := x"55E"; 
		s_E689_C1_L				  :std_logic_vector(11 downto 0) := x"560"; 
		s_E690_C1_L				  :std_logic_vector(11 downto 0) := x"562"; 
		s_E691_C1_L				  :std_logic_vector(11 downto 0) := x"564"; 
		s_E692_C1_L				  :std_logic_vector(11 downto 0) := x"566"; 
		s_E693_C1_L				  :std_logic_vector(11 downto 0) := x"568"; 
		s_E694_C1_L				  :std_logic_vector(11 downto 0) := x"56A"; 
		s_E695_C1_L				  :std_logic_vector(11 downto 0) := x"56C"; 
		s_E696_C1_L				  :std_logic_vector(11 downto 0) := x"56E"; 
		s_E697_C1_L				  :std_logic_vector(11 downto 0) := x"570"; 
		s_E698_C1_L				  :std_logic_vector(11 downto 0) := x"572"; 
		s_E699_C1_L				  :std_logic_vector(11 downto 0) := x"574"; 
		s_E700_C1_L				  :std_logic_vector(11 downto 0) := x"576"; 
		s_E701_C1_L				  :std_logic_vector(11 downto 0) := x"578"; 
		s_E702_C1_L				  :std_logic_vector(11 downto 0) := x"57A"; 
		s_E703_C1_L				  :std_logic_vector(11 downto 0) := x"57C"; 
		s_E704_C1_L				  :std_logic_vector(11 downto 0) := x"57E"; 
		s_E705_C1_L				  :std_logic_vector(11 downto 0) := x"580"; 
		s_E706_C1_L				  :std_logic_vector(11 downto 0) := x"582"; 
		s_E707_C1_L				  :std_logic_vector(11 downto 0) := x"584"; 
		s_E708_C1_L				  :std_logic_vector(11 downto 0) := x"586"; 
		s_E709_C1_L				  :std_logic_vector(11 downto 0) := x"588"; 
		s_E710_C1_L				  :std_logic_vector(11 downto 0) := x"58A"; 
		s_E711_C1_L				  :std_logic_vector(11 downto 0) := x"58C"; 
		s_E712_C1_L				  :std_logic_vector(11 downto 0) := x"58E"; 
		s_E713_C1_L				  :std_logic_vector(11 downto 0) := x"590"; 
		s_E714_C1_L				  :std_logic_vector(11 downto 0) := x"592"; 
		s_E715_C1_L				  :std_logic_vector(11 downto 0) := x"594"; 
		s_E716_C1_L				  :std_logic_vector(11 downto 0) := x"596"; 
		s_E717_C1_L				  :std_logic_vector(11 downto 0) := x"598"; 
		s_E718_C1_L				  :std_logic_vector(11 downto 0) := x"59A"; 
		s_E719_C1_L				  :std_logic_vector(11 downto 0) := x"59C"; 
		s_E720_C1_L				  :std_logic_vector(11 downto 0) := x"59E"; 
		s_E721_C1_L				  :std_logic_vector(11 downto 0) := x"5A0"; 
		s_E722_C1_L				  :std_logic_vector(11 downto 0) := x"5A2"; 
		s_E723_C1_L				  :std_logic_vector(11 downto 0) := x"5A4"; 
		s_E724_C1_L				  :std_logic_vector(11 downto 0) := x"5A6"; 
		s_E725_C1_L				  :std_logic_vector(11 downto 0) := x"5A8"; 
		s_E726_C1_L				  :std_logic_vector(11 downto 0) := x"5AA"; 
		s_E727_C1_L				  :std_logic_vector(11 downto 0) := x"5AC"; 
		s_E728_C1_L				  :std_logic_vector(11 downto 0) := x"5AE"; 
		s_E729_C1_L				  :std_logic_vector(11 downto 0) := x"5B0"; 
		s_E730_C1_L				  :std_logic_vector(11 downto 0) := x"5B2"; 
		s_E731_C1_L				  :std_logic_vector(11 downto 0) := x"5B4"; 
		s_E732_C1_L				  :std_logic_vector(11 downto 0) := x"5B6"; 
		s_E733_C1_L				  :std_logic_vector(11 downto 0) := x"5B8"; 
		s_E734_C1_L				  :std_logic_vector(11 downto 0) := x"5BA"; 
		s_E735_C1_L				  :std_logic_vector(11 downto 0) := x"5BC"; 
		s_E736_C1_L				  :std_logic_vector(11 downto 0) := x"5BE"; 
		s_E737_C1_L				  :std_logic_vector(11 downto 0) := x"5C0"; 
		s_E738_C1_L				  :std_logic_vector(11 downto 0) := x"5C2"; 
		s_E739_C1_L				  :std_logic_vector(11 downto 0) := x"5C4"; 
		s_E740_C1_L				  :std_logic_vector(11 downto 0) := x"5C6"; 
		s_E741_C1_L				  :std_logic_vector(11 downto 0) := x"5C8"; 
		s_E742_C1_L				  :std_logic_vector(11 downto 0) := x"5CA"; 
		s_E743_C1_L				  :std_logic_vector(11 downto 0) := x"5CC"; 
		s_E744_C1_L				  :std_logic_vector(11 downto 0) := x"5CE"; 
		s_E745_C1_L				  :std_logic_vector(11 downto 0) := x"5D0"; 
		s_E746_C1_L				  :std_logic_vector(11 downto 0) := x"5D2"; 
		s_E747_C1_L				  :std_logic_vector(11 downto 0) := x"5D4"; 
		s_E748_C1_L				  :std_logic_vector(11 downto 0) := x"5D6"; 
		s_E749_C1_L				  :std_logic_vector(11 downto 0) := x"5D8"; 
		s_E750_C1_L				  :std_logic_vector(11 downto 0) := x"5DA"; 
		s_E751_C1_L				  :std_logic_vector(11 downto 0) := x"5DC"; 
		s_E752_C1_L				  :std_logic_vector(11 downto 0) := x"5DE"; 
		s_E753_C1_L				  :std_logic_vector(11 downto 0) := x"5E0"; 
		s_E754_C1_L				  :std_logic_vector(11 downto 0) := x"5E2"; 
		s_E755_C1_L				  :std_logic_vector(11 downto 0) := x"5E4"; 
		s_E756_C1_L				  :std_logic_vector(11 downto 0) := x"5E6"; 
		s_E757_C1_L				  :std_logic_vector(11 downto 0) := x"5E8"; 
		s_E758_C1_L				  :std_logic_vector(11 downto 0) := x"5EA"; 
		s_E759_C1_L				  :std_logic_vector(11 downto 0) := x"5EC"; 
		s_E760_C1_L				  :std_logic_vector(11 downto 0) := x"5EE"; 
		s_E761_C1_L				  :std_logic_vector(11 downto 0) := x"5F0"; 
		s_E762_C1_L				  :std_logic_vector(11 downto 0) := x"5F2"; 
		s_E763_C1_L				  :std_logic_vector(11 downto 0) := x"5F4"; 
		s_E764_C1_L				  :std_logic_vector(11 downto 0) := x"5F6"; 
		s_E765_C1_L				  :std_logic_vector(11 downto 0) := x"5F8"; 
		s_E766_C1_L				  :std_logic_vector(11 downto 0) := x"5FA"; 
		s_E767_C1_L				  :std_logic_vector(11 downto 0) := x"5FC"; 
		s_E768_C1_L				  :std_logic_vector(11 downto 0) := x"5FE"; 
		s_E769_C1_L				  :std_logic_vector(11 downto 0) := x"600"; 
		s_E770_C1_L				  :std_logic_vector(11 downto 0) := x"602"; 
		s_E771_C1_L				  :std_logic_vector(11 downto 0) := x"604"; 
		s_E772_C1_L				  :std_logic_vector(11 downto 0) := x"606"; 
		s_E773_C1_L				  :std_logic_vector(11 downto 0) := x"608"; 
		s_E774_C1_L				  :std_logic_vector(11 downto 0) := x"60A"; 
		s_E775_C1_L				  :std_logic_vector(11 downto 0) := x"60C"; 
		s_E776_C1_L				  :std_logic_vector(11 downto 0) := x"60E"; 
		s_E777_C1_L				  :std_logic_vector(11 downto 0) := x"610"; 
		s_E778_C1_L				  :std_logic_vector(11 downto 0) := x"612"; 
		s_E779_C1_L				  :std_logic_vector(11 downto 0) := x"614"; 
		s_E780_C1_L				  :std_logic_vector(11 downto 0) := x"616"; 
		s_E781_C1_L				  :std_logic_vector(11 downto 0) := x"618"; 
		s_E782_C1_L				  :std_logic_vector(11 downto 0) := x"61A"; 
		s_E783_C1_L				  :std_logic_vector(11 downto 0) := x"61C"; 
		s_E784_C1_L				  :std_logic_vector(11 downto 0) := x"61E"; 
		s_E785_C1_L				  :std_logic_vector(11 downto 0) := x"620"; 
		s_E786_C1_L				  :std_logic_vector(11 downto 0) := x"622"; 
		s_E787_C1_L				  :std_logic_vector(11 downto 0) := x"624"; 
		s_E788_C1_L				  :std_logic_vector(11 downto 0) := x"626"; 
		s_E789_C1_L				  :std_logic_vector(11 downto 0) := x"628"; 
		s_E790_C1_L				  :std_logic_vector(11 downto 0) := x"62A"; 
		s_E791_C1_L				  :std_logic_vector(11 downto 0) := x"62C"; 
		s_E792_C1_L				  :std_logic_vector(11 downto 0) := x"62E"; 
		s_E793_C1_L				  :std_logic_vector(11 downto 0) := x"630"; 
		s_E794_C1_L				  :std_logic_vector(11 downto 0) := x"632"; 
		s_E795_C1_L				  :std_logic_vector(11 downto 0) := x"634"; 
		s_E796_C1_L				  :std_logic_vector(11 downto 0) := x"636"; 
		s_E797_C1_L				  :std_logic_vector(11 downto 0) := x"638"; 
		s_E798_C1_L				  :std_logic_vector(11 downto 0) := x"63A"; 
		s_E799_C1_L				  :std_logic_vector(11 downto 0) := x"63C"; 
		s_E800_C1_L				  :std_logic_vector(11 downto 0) := x"63E"; 
		s_E801_C1_L				  :std_logic_vector(11 downto 0) := x"640"; 
		s_E802_C1_L				  :std_logic_vector(11 downto 0) := x"642"; 
		s_E803_C1_L				  :std_logic_vector(11 downto 0) := x"644"; 
		s_E804_C1_L				  :std_logic_vector(11 downto 0) := x"646"; 
		s_E805_C1_L				  :std_logic_vector(11 downto 0) := x"648"; 
		s_E806_C1_L				  :std_logic_vector(11 downto 0) := x"64A"; 
		s_E807_C1_L				  :std_logic_vector(11 downto 0) := x"64C"; 
		s_E808_C1_L				  :std_logic_vector(11 downto 0) := x"64E"; 
		s_E809_C1_L				  :std_logic_vector(11 downto 0) := x"650"; 
		s_E810_C1_L				  :std_logic_vector(11 downto 0) := x"652"; 
		s_E811_C1_L				  :std_logic_vector(11 downto 0) := x"654"; 
		s_E812_C1_L				  :std_logic_vector(11 downto 0) := x"656"; 
		s_E813_C1_L				  :std_logic_vector(11 downto 0) := x"658"; 
		s_E814_C1_L				  :std_logic_vector(11 downto 0) := x"65A"; 
		s_E815_C1_L				  :std_logic_vector(11 downto 0) := x"65C"; 
		s_E816_C1_L				  :std_logic_vector(11 downto 0) := x"65E"; 
		s_E817_C1_L				  :std_logic_vector(11 downto 0) := x"660"; 
		s_E818_C1_L				  :std_logic_vector(11 downto 0) := x"662"; 
		s_E819_C1_L				  :std_logic_vector(11 downto 0) := x"664"; 
		s_E820_C1_L				  :std_logic_vector(11 downto 0) := x"666"; 
		s_E821_C1_L				  :std_logic_vector(11 downto 0) := x"668"; 
		s_E822_C1_L				  :std_logic_vector(11 downto 0) := x"66A"; 
		s_E823_C1_L				  :std_logic_vector(11 downto 0) := x"66C"; 
		s_E824_C1_L				  :std_logic_vector(11 downto 0) := x"66E"; 
		s_E825_C1_L				  :std_logic_vector(11 downto 0) := x"670"; 
		s_E826_C1_L				  :std_logic_vector(11 downto 0) := x"672"; 
		s_E827_C1_L				  :std_logic_vector(11 downto 0) := x"674"; 
		s_E828_C1_L				  :std_logic_vector(11 downto 0) := x"676"; 
		s_E829_C1_L				  :std_logic_vector(11 downto 0) := x"678"; 
		s_E830_C1_L				  :std_logic_vector(11 downto 0) := x"67A"; 
		s_E831_C1_L				  :std_logic_vector(11 downto 0) := x"67C"; 
		s_E832_C1_L				  :std_logic_vector(11 downto 0) := x"67E"; 
		s_E833_C1_L				  :std_logic_vector(11 downto 0) := x"680"; 
		s_E834_C1_L				  :std_logic_vector(11 downto 0) := x"682"; 
		s_E835_C1_L				  :std_logic_vector(11 downto 0) := x"684"; 
		s_E836_C1_L				  :std_logic_vector(11 downto 0) := x"686"; 
		s_E837_C1_L				  :std_logic_vector(11 downto 0) := x"688"; 
		s_E838_C1_L				  :std_logic_vector(11 downto 0) := x"68A"; 
		s_E839_C1_L				  :std_logic_vector(11 downto 0) := x"68C"; 
		s_E840_C1_L				  :std_logic_vector(11 downto 0) := x"68E"; 
		s_E841_C1_L				  :std_logic_vector(11 downto 0) := x"690"; 
		s_E842_C1_L				  :std_logic_vector(11 downto 0) := x"692"; 
		s_E843_C1_L				  :std_logic_vector(11 downto 0) := x"694"; 
		s_E844_C1_L				  :std_logic_vector(11 downto 0) := x"696"; 
		s_E845_C1_L				  :std_logic_vector(11 downto 0) := x"698"; 
		s_E846_C1_L				  :std_logic_vector(11 downto 0) := x"69A"; 
		s_E847_C1_L				  :std_logic_vector(11 downto 0) := x"69C"; 
		s_E848_C1_L				  :std_logic_vector(11 downto 0) := x"69E"; 
		s_E849_C1_L				  :std_logic_vector(11 downto 0) := x"6A0"; 
		s_E850_C1_L				  :std_logic_vector(11 downto 0) := x"6A2"; 
		s_E851_C1_L				  :std_logic_vector(11 downto 0) := x"6A4"; 
		s_E852_C1_L				  :std_logic_vector(11 downto 0) := x"6A6"; 
		s_E853_C1_L				  :std_logic_vector(11 downto 0) := x"6A8"; 
		s_E854_C1_L				  :std_logic_vector(11 downto 0) := x"6AA"; 
		s_E855_C1_L				  :std_logic_vector(11 downto 0) := x"6AC"; 
		s_E856_C1_L				  :std_logic_vector(11 downto 0) := x"6AE"; 
		s_E857_C1_L				  :std_logic_vector(11 downto 0) := x"6B0"; 
		s_E858_C1_L				  :std_logic_vector(11 downto 0) := x"6B2"; 
		s_E859_C1_L				  :std_logic_vector(11 downto 0) := x"6B4"; 
		s_E860_C1_L				  :std_logic_vector(11 downto 0) := x"6B6"; 
		s_E861_C1_L				  :std_logic_vector(11 downto 0) := x"6B8"; 
		s_E862_C1_L				  :std_logic_vector(11 downto 0) := x"6BA"; 
		s_E863_C1_L				  :std_logic_vector(11 downto 0) := x"6BC"; 
		s_E864_C1_L				  :std_logic_vector(11 downto 0) := x"6BE"; 
		s_E865_C1_L				  :std_logic_vector(11 downto 0) := x"6C0"; 
		s_E866_C1_L				  :std_logic_vector(11 downto 0) := x"6C2"; 
		s_E867_C1_L				  :std_logic_vector(11 downto 0) := x"6C4"; 
		s_E868_C1_L				  :std_logic_vector(11 downto 0) := x"6C6"; 
		s_E869_C1_L				  :std_logic_vector(11 downto 0) := x"6C8"; 
		s_E870_C1_L				  :std_logic_vector(11 downto 0) := x"6CA"; 
		s_E871_C1_L				  :std_logic_vector(11 downto 0) := x"6CC"; 
		s_E872_C1_L				  :std_logic_vector(11 downto 0) := x"6CE"; 
		s_E873_C1_L				  :std_logic_vector(11 downto 0) := x"6D0"; 
		s_E874_C1_L				  :std_logic_vector(11 downto 0) := x"6D2"; 
		s_E875_C1_L				  :std_logic_vector(11 downto 0) := x"6D4"; 
		s_E876_C1_L				  :std_logic_vector(11 downto 0) := x"6D6"; 
		s_E877_C1_L				  :std_logic_vector(11 downto 0) := x"6D8"; 
		s_E878_C1_L				  :std_logic_vector(11 downto 0) := x"6DA"; 
		s_E879_C1_L				  :std_logic_vector(11 downto 0) := x"6DC"; 
		s_E880_C1_L				  :std_logic_vector(11 downto 0) := x"6DE"; 
		s_E881_C1_L				  :std_logic_vector(11 downto 0) := x"6E0"; 
		s_E882_C1_L				  :std_logic_vector(11 downto 0) := x"6E2"; 
		s_E883_C1_L				  :std_logic_vector(11 downto 0) := x"6E4"; 
		s_E884_C1_L				  :std_logic_vector(11 downto 0) := x"6E6"; 
		s_E885_C1_L				  :std_logic_vector(11 downto 0) := x"6E8"; 
		s_E886_C1_L				  :std_logic_vector(11 downto 0) := x"6EA"; 
		s_E887_C1_L				  :std_logic_vector(11 downto 0) := x"6EC"; 
		s_E888_C1_L				  :std_logic_vector(11 downto 0) := x"6EE"; 
		s_E889_C1_L				  :std_logic_vector(11 downto 0) := x"6F0"; 
		s_E890_C1_L				  :std_logic_vector(11 downto 0) := x"6F2"; 
		s_E891_C1_L				  :std_logic_vector(11 downto 0) := x"6F4"; 
		s_E892_C1_L				  :std_logic_vector(11 downto 0) := x"6F6"; 
		s_E893_C1_L				  :std_logic_vector(11 downto 0) := x"6F8"; 
		s_E894_C1_L				  :std_logic_vector(11 downto 0) := x"6FA"; 
		s_E895_C1_L				  :std_logic_vector(11 downto 0) := x"6FC"; 
		s_E896_C1_L				  :std_logic_vector(11 downto 0) := x"6FE"; 
		s_E897_C1_L				  :std_logic_vector(11 downto 0) := x"700"; 
		s_E898_C1_L				  :std_logic_vector(11 downto 0) := x"702"; 
		s_E899_C1_L				  :std_logic_vector(11 downto 0) := x"704"; 
		s_E900_C1_L				  :std_logic_vector(11 downto 0) := x"706"; 
		s_E901_C1_L				  :std_logic_vector(11 downto 0) := x"708"; 
		s_E902_C1_L				  :std_logic_vector(11 downto 0) := x"70A"; 
		s_E903_C1_L				  :std_logic_vector(11 downto 0) := x"70C"; 
		s_E904_C1_L				  :std_logic_vector(11 downto 0) := x"70E"; 
		s_E905_C1_L				  :std_logic_vector(11 downto 0) := x"710"; 
		s_E906_C1_L				  :std_logic_vector(11 downto 0) := x"712"; 
		s_E907_C1_L				  :std_logic_vector(11 downto 0) := x"714"; 
		s_E908_C1_L				  :std_logic_vector(11 downto 0) := x"716"; 
		s_E909_C1_L				  :std_logic_vector(11 downto 0) := x"718"; 
		s_E910_C1_L				  :std_logic_vector(11 downto 0) := x"71A"; 
		s_E911_C1_L				  :std_logic_vector(11 downto 0) := x"71C"; 
		s_E912_C1_L				  :std_logic_vector(11 downto 0) := x"71E"; 
		s_E913_C1_L				  :std_logic_vector(11 downto 0) := x"720"; 
		s_E914_C1_L				  :std_logic_vector(11 downto 0) := x"722"; 
		s_E915_C1_L				  :std_logic_vector(11 downto 0) := x"724"; 
		s_E916_C1_L				  :std_logic_vector(11 downto 0) := x"726"; 
		s_E917_C1_L				  :std_logic_vector(11 downto 0) := x"728"; 
		s_E918_C1_L				  :std_logic_vector(11 downto 0) := x"72A"; 
		s_E919_C1_L				  :std_logic_vector(11 downto 0) := x"72C"; 
		s_E920_C1_L				  :std_logic_vector(11 downto 0) := x"72E"; 
		s_E921_C1_L				  :std_logic_vector(11 downto 0) := x"730"; 
		s_E922_C1_L				  :std_logic_vector(11 downto 0) := x"732"; 
		s_E923_C1_L				  :std_logic_vector(11 downto 0) := x"734"; 
		s_E924_C1_L				  :std_logic_vector(11 downto 0) := x"736"; 
		s_E925_C1_L				  :std_logic_vector(11 downto 0) := x"738"; 
		s_E926_C1_L				  :std_logic_vector(11 downto 0) := x"73A"; 
		s_E927_C1_L				  :std_logic_vector(11 downto 0) := x"73C"; 
		s_E928_C1_L				  :std_logic_vector(11 downto 0) := x"73E"; 
		s_E929_C1_L				  :std_logic_vector(11 downto 0) := x"740"; 
		s_E930_C1_L				  :std_logic_vector(11 downto 0) := x"742"; 
		s_E931_C1_L				  :std_logic_vector(11 downto 0) := x"744"; 
		s_E932_C1_L				  :std_logic_vector(11 downto 0) := x"746"; 
		s_E933_C1_L				  :std_logic_vector(11 downto 0) := x"748"; 
		s_E934_C1_L				  :std_logic_vector(11 downto 0) := x"74A"; 
		s_E935_C1_L				  :std_logic_vector(11 downto 0) := x"74C"; 
		s_E936_C1_L				  :std_logic_vector(11 downto 0) := x"74E"; 
		s_E937_C1_L				  :std_logic_vector(11 downto 0) := x"750"; 
		s_E938_C1_L				  :std_logic_vector(11 downto 0) := x"752"; 
		s_E939_C1_L				  :std_logic_vector(11 downto 0) := x"754"; 
		s_E940_C1_L				  :std_logic_vector(11 downto 0) := x"756"; 
		s_E941_C1_L				  :std_logic_vector(11 downto 0) := x"758"; 
		s_E942_C1_L				  :std_logic_vector(11 downto 0) := x"75A"; 
		s_E943_C1_L				  :std_logic_vector(11 downto 0) := x"75C"; 
		s_E944_C1_L				  :std_logic_vector(11 downto 0) := x"75E"; 
		s_E945_C1_L				  :std_logic_vector(11 downto 0) := x"760"; 
		s_E946_C1_L				  :std_logic_vector(11 downto 0) := x"762"; 
		s_E947_C1_L				  :std_logic_vector(11 downto 0) := x"764"; 
		s_E948_C1_L				  :std_logic_vector(11 downto 0) := x"766"; 
		s_E949_C1_L				  :std_logic_vector(11 downto 0) := x"768"; 
		s_E950_C1_L				  :std_logic_vector(11 downto 0) := x"76A"; 
		s_E951_C1_L				  :std_logic_vector(11 downto 0) := x"76C"; 
		s_E952_C1_L				  :std_logic_vector(11 downto 0) := x"76E"; 
		s_E953_C1_L				  :std_logic_vector(11 downto 0) := x"770"; 
		s_E954_C1_L				  :std_logic_vector(11 downto 0) := x"772"; 
		s_E955_C1_L				  :std_logic_vector(11 downto 0) := x"774"; 
		s_E956_C1_L				  :std_logic_vector(11 downto 0) := x"776"; 
		s_E957_C1_L				  :std_logic_vector(11 downto 0) := x"778"; 
		s_E958_C1_L				  :std_logic_vector(11 downto 0) := x"77A"; 
		s_E959_C1_L				  :std_logic_vector(11 downto 0) := x"77C"; 
		s_E960_C1_L				  :std_logic_vector(11 downto 0) := x"77E"; 
		s_E961_C1_L				  :std_logic_vector(11 downto 0) := x"780"; 
		s_E962_C1_L				  :std_logic_vector(11 downto 0) := x"782"; 
		s_E963_C1_L				  :std_logic_vector(11 downto 0) := x"784"; 
		s_E964_C1_L				  :std_logic_vector(11 downto 0) := x"786"; 
		s_E965_C1_L				  :std_logic_vector(11 downto 0) := x"788"; 
		s_E966_C1_L				  :std_logic_vector(11 downto 0) := x"78A"; 
		s_E967_C1_L				  :std_logic_vector(11 downto 0) := x"78C"; 
		s_E968_C1_L				  :std_logic_vector(11 downto 0) := x"78E"; 
		s_E969_C1_L				  :std_logic_vector(11 downto 0) := x"790"; 
		s_E970_C1_L				  :std_logic_vector(11 downto 0) := x"792"; 
		s_E971_C1_L				  :std_logic_vector(11 downto 0) := x"794"; 
		s_E972_C1_L				  :std_logic_vector(11 downto 0) := x"796"; 
		s_E973_C1_L				  :std_logic_vector(11 downto 0) := x"798"; 
		s_E974_C1_L				  :std_logic_vector(11 downto 0) := x"79A"; 
		s_E975_C1_L				  :std_logic_vector(11 downto 0) := x"79C"; 
		s_E976_C1_L				  :std_logic_vector(11 downto 0) := x"79E"; 
		s_E977_C1_L				  :std_logic_vector(11 downto 0) := x"7A0"; 
		s_E978_C1_L				  :std_logic_vector(11 downto 0) := x"7A2"; 
		s_E979_C1_L				  :std_logic_vector(11 downto 0) := x"7A4"; 
		s_E980_C1_L				  :std_logic_vector(11 downto 0) := x"7A6"; 
		s_E981_C1_L				  :std_logic_vector(11 downto 0) := x"7A8"; 
		s_E982_C1_L				  :std_logic_vector(11 downto 0) := x"7AA"; 
		s_E983_C1_L				  :std_logic_vector(11 downto 0) := x"7AC"; 
		s_E984_C1_L				  :std_logic_vector(11 downto 0) := x"7AE"; 
		s_E985_C1_L				  :std_logic_vector(11 downto 0) := x"7B0"; 
		s_E986_C1_L				  :std_logic_vector(11 downto 0) := x"7B2"; 
		s_E987_C1_L				  :std_logic_vector(11 downto 0) := x"7B4"; 
		s_E988_C1_L				  :std_logic_vector(11 downto 0) := x"7B6"; 
		s_E989_C1_L				  :std_logic_vector(11 downto 0) := x"7B8"; 
		s_E990_C1_L				  :std_logic_vector(11 downto 0) := x"7BA"; 
		s_E991_C1_L				  :std_logic_vector(11 downto 0) := x"7BC"; 
		s_E992_C1_L				  :std_logic_vector(11 downto 0) := x"7BE"; 
		s_E993_C1_L				  :std_logic_vector(11 downto 0) := x"7C0"; 
		s_E994_C1_L				  :std_logic_vector(11 downto 0) := x"7C2"; 
		s_E995_C1_L				  :std_logic_vector(11 downto 0) := x"7C4"; 
		s_E996_C1_L				  :std_logic_vector(11 downto 0) := x"7C6"; 
		s_E997_C1_L				  :std_logic_vector(11 downto 0) := x"7C8"; 
		s_E998_C1_L				  :std_logic_vector(11 downto 0) := x"7CA"; 
		s_E999_C1_L				  :std_logic_vector(11 downto 0) := x"7CC"; 
		s_E1000_C1_L			  :std_logic_vector(11 downto 0) := x"7CE"; 
		s_E1001_C1_L			  :std_logic_vector(11 downto 0) := x"7D0"; 
		s_E1002_C1_L			  :std_logic_vector(11 downto 0) := x"7D2"; 
		s_E1003_C1_L			  :std_logic_vector(11 downto 0) := x"7D4"; 
		s_E1004_C1_L			  :std_logic_vector(11 downto 0) := x"7D6"; 
		s_E1005_C1_L			  :std_logic_vector(11 downto 0) := x"7D8"; 
		s_E1006_C1_L			  :std_logic_vector(11 downto 0) := x"7DA"; 
		s_E1007_C1_L			  :std_logic_vector(11 downto 0) := x"7DC"; 
		s_E1008_C1_L			  :std_logic_vector(11 downto 0) := x"7DE"; 
		s_E1009_C1_L			  :std_logic_vector(11 downto 0) := x"7E0"; 
		s_E1010_C1_L			  :std_logic_vector(11 downto 0) := x"7E2"; 
		s_E1011_C1_L			  :std_logic_vector(11 downto 0) := x"7E4"; 
		s_E1012_C1_L			  :std_logic_vector(11 downto 0) := x"7E6"; 
		s_E1013_C1_L			  :std_logic_vector(11 downto 0) := x"7E8"; 
		s_E1014_C1_L			  :std_logic_vector(11 downto 0) := x"7EA"; 
		s_E1015_C1_L			  :std_logic_vector(11 downto 0) := x"7EC"; 
		s_E1016_C1_L			  :std_logic_vector(11 downto 0) := x"7EE"; 
		s_E1017_C1_L			  :std_logic_vector(11 downto 0) := x"7F0"; 
		s_E1018_C1_L			  :std_logic_vector(11 downto 0) := x"7F2"; 
		s_E1019_C1_L			  :std_logic_vector(11 downto 0) := x"7F4"; 
		s_E1020_C1_L			  :std_logic_vector(11 downto 0) := x"7F6"; 
		s_E1021_C1_L			  :std_logic_vector(11 downto 0) := x"7F8"; 
		s_E1022_C1_L			  :std_logic_vector(11 downto 0) := x"7FA"; 
		s_E1023_C1_L			  :std_logic_vector(11 downto 0) := x"7FC"; 
		s_E1024_C1_L			  :std_logic_vector(11 downto 0) := x"7FE"; 
                                                                    
		s_E1_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"7FF";
		s_E1_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"801";
		s_E2_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"803";
		s_E3_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"805";
		s_E4_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"807";
		s_E5_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"809";
		s_E6_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"80B";
		s_E7_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"80D";
		s_E8_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"80F";
		s_E9_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"811";
		s_E10_C1_H_Pos       	  :std_logic_vector(11 downto 0) := x"813";
		s_E11_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"815";
		s_E12_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"817";
		s_E13_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"819";
		s_E14_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"81B";
		s_E15_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"81D";
		s_E16_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"81F";
		s_E17_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"821";
		s_E18_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"823";
		s_E19_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"825";
		s_E20_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"827";
		s_E21_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"829";
		s_E22_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"82B";
		s_E23_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"82D";
		s_E24_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"82F";
		s_E25_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"831";
		s_E26_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"833";
		s_E27_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"835";
		s_E28_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"837";
		s_E29_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"839";
		s_E30_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"83B";
		s_E31_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"83D";
		s_E32_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"83F";
		s_E33_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"841";
		s_E34_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"843";
		s_E35_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"845";
		s_E36_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"847";
		s_E37_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"849";
		s_E38_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"84B";
		s_E39_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"84D";
		s_E40_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"84F";
		s_E41_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"851";
		s_E42_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"853";
		s_E43_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"855";
		s_E44_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"857";
		s_E45_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"859";
		s_E46_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"85B";
		s_E47_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"85D";
		s_E48_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"85F";
		s_E49_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"861";
		s_E50_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"863";
		s_E51_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"865";
		s_E52_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"867";
		s_E53_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"869";
		s_E54_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"86B";
		s_E55_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"86D";
		s_E56_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"86F";
		s_E57_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"871";
		s_E58_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"873";
		s_E59_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"875";
		s_E60_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"877";
		s_E61_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"879";
		s_E62_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"87B";
		s_E63_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"87D";
		s_E64_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"87F";
		s_E65_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"881";
		s_E66_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"883";
		s_E67_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"885";
		s_E68_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"887";
		s_E69_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"889";
		s_E70_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"88B";
		s_E71_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"88D";
		s_E72_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"88F";
		s_E73_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"891";
		s_E74_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"893";
		s_E75_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"895";
		s_E76_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"897";
		s_E77_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"899";
		s_E78_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"89B";
		s_E79_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"89D";
		s_E80_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"89F";
		s_E81_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8A1";
		s_E82_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8A3";
		s_E83_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8A5";
		s_E84_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8A7";
		s_E85_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8A9";
		s_E86_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8AB";
		s_E87_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8AD";
		s_E88_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8AF";
		s_E89_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8B1";
		s_E90_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8B3";
		s_E91_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8B5";
		s_E92_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8B7";
		s_E93_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8B9";
		s_E94_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8BB";
		s_E95_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8BD";
		s_E96_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8BF";
		s_E97_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8C1";
		s_E98_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8C3";
		s_E99_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8C5";
		s_E100_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8C7";
		s_E101_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8C9";
		s_E102_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8CB";
		s_E103_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8CD";
		s_E104_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8CF";
		s_E105_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8D1";
		s_E106_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8D3";
		s_E107_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8D5";
		s_E108_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8D7";
		s_E109_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8D9";
		s_E110_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8DB";
		s_E111_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8DD";
		s_E112_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8DF";
		s_E113_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8E1";
		s_E114_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8E3";
		s_E115_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8E5";
		s_E116_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8E7";
		s_E117_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8E9";
		s_E118_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8EB";
		s_E119_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8ED";
		s_E120_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8EF";
		s_E121_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8F1";
		s_E122_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8F3";
		s_E123_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8F5";
		s_E124_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8F7";
		s_E125_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8F9";
		s_E126_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8FB";
		s_E127_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8FD";
		s_E128_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8FF";
		s_E129_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"901";
		s_E130_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"903";
		s_E131_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"905";
		s_E132_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"907";
		s_E133_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"909";
		s_E134_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"90B";
		s_E135_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"90D";
		s_E136_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"90F";
		s_E137_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"911";
		s_E138_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"913";
		s_E139_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"915";
		s_E140_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"917";
		s_E141_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"919";
		s_E142_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"91B";
		s_E143_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"91D";
		s_E144_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"91F";
		s_E145_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"921";
		s_E146_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"923";
		s_E147_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"925";
		s_E148_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"927";
		s_E149_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"929";
		s_E150_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"92B";
		s_E151_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"92D";
		s_E152_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"92F";
		s_E153_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"931";
		s_E154_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"933";
		s_E155_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"935";
		s_E156_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"937";
		s_E157_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"939";
		s_E158_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"93B";
		s_E159_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"93D";
		s_E160_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"93F";
		s_E161_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"941";
		s_E162_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"943";
		s_E163_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"945";
		s_E164_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"947";
		s_E165_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"949";
		s_E166_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"94B";
		s_E167_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"94D";
		s_E168_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"94F";
		s_E169_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"951";
		s_E170_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"953";
		s_E171_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"955";
		s_E172_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"957";
		s_E173_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"959";
		s_E174_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"95B";
		s_E175_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"95D";
		s_E176_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"95F";
		s_E177_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"961";
		s_E178_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"963";
		s_E179_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"965";
		s_E180_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"967";
		s_E181_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"969";
		s_E182_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"96B";
		s_E183_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"96D";
		s_E184_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"96F";
		s_E185_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"971";
		s_E186_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"973";
		s_E187_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"975";
		s_E188_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"977";
		s_E189_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"979";
		s_E190_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"97B";
		s_E191_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"97D";
		s_E192_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"97F";
		s_E193_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"981";
		s_E194_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"983";
		s_E195_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"985";
		s_E196_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"987";
		s_E197_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"989";
		s_E198_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"98B";
		s_E199_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"98D";
		s_E200_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"98F";
		s_E201_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"991";
		s_E202_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"993";
		s_E203_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"995";
		s_E204_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"997";
		s_E205_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"999";
		s_E206_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"99B";
		s_E207_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"99D";
		s_E208_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"99F";
		s_E209_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9A1";
		s_E210_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9A3";
		s_E211_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9A5";
		s_E212_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9A7";
		s_E213_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9A9";
		s_E214_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9AB";
		s_E215_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9AD";
		s_E216_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9AF";
		s_E217_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9B1";
		s_E218_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9B3";
		s_E219_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9B5";
		s_E220_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9B7";
		s_E221_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9B9";
		s_E222_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9BB";
		s_E223_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9BD";
		s_E224_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9BF";
		s_E225_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9C1";
		s_E226_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9C3";
		s_E227_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9C5";
		s_E228_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9C7";
		s_E229_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9C9";
		s_E230_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9CB";
		s_E231_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9CD";
		s_E232_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9CF";
		s_E233_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9D1";
		s_E234_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9D3";
		s_E235_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9D5";
		s_E236_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9D7";
		s_E237_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9D9";
		s_E238_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9DB";
		s_E239_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9DD";
		s_E240_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9DF";
		s_E241_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9E1";
		s_E242_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9E3";
		s_E243_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9E5";
		s_E244_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9E7";
		s_E245_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9E9";
		s_E246_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9EB";
		s_E247_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9ED";
		s_E248_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9EF";
		s_E249_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9F1";
		s_E250_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9F3";
		s_E251_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9F5";
		s_E252_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9F7";
		s_E253_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9F9";
		s_E254_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9FB";
		s_E255_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9FD";
		s_E256_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9FF";
		s_E257_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A01";
		s_E258_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A03";
		s_E259_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A05";
		s_E260_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A07";
		s_E261_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A09";
		s_E262_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A0B";
		s_E263_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A0D";
		s_E264_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A0F";
		s_E265_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A11";
		s_E266_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A13";
		s_E267_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A15";
		s_E268_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A17";
		s_E269_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A19";
		s_E270_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A1B";
		s_E271_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A1D";
		s_E272_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A1F";
		s_E273_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A21";
		s_E274_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A23";
		s_E275_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A25";
		s_E276_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A27";
		s_E277_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A29";
		s_E278_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A2B";
		s_E279_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A2D";
		s_E280_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A2F";
		s_E281_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A31";
		s_E282_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A33";
		s_E283_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A35";
		s_E284_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A37";
		s_E285_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A39";
		s_E286_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A3B";
		s_E287_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A3D";
		s_E288_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A3F";
		s_E289_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A41";
		s_E290_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A43";
		s_E291_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A45";
		s_E292_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A47";
		s_E293_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A49";
		s_E294_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A4B";
		s_E295_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A4D";
		s_E296_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A4F";
		s_E297_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A51";
		s_E298_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A53";
		s_E299_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A55";
		s_E300_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A57";
		s_E301_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A59";
		s_E302_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A5B";
		s_E303_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A5D";
		s_E304_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A5F";
		s_E305_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A61";
		s_E306_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A63";
		s_E307_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A65";
		s_E308_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A67";
		s_E309_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A69";
		s_E310_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A6B";
		s_E311_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A6D";
		s_E312_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A6F";
		s_E313_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A71";
		s_E314_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A73";
		s_E315_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A75";
		s_E316_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A77";
		s_E317_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A79";
		s_E318_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A7B";
		s_E319_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A7D";
		s_E320_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A7F";
		s_E321_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A81";
		s_E322_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A83";
		s_E323_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A85";
		s_E324_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A87";
		s_E325_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A89";
		s_E326_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A8B";
		s_E327_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A8D";
		s_E328_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A8F";
		s_E329_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A91";
		s_E330_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A93";
		s_E331_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A95";
		s_E332_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A97";
		s_E333_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A99";
		s_E334_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A9B";
		s_E335_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A9D";
		s_E336_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A9F";
		s_E337_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AA1";
		s_E338_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AA3";
		s_E339_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AA5";
		s_E340_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AA7";
		s_E341_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AA9";
		s_E342_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AAB";
		s_E343_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AAD";
		s_E344_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AAF";
		s_E345_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AB1";
		s_E346_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AB3";
		s_E347_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AB5";
		s_E348_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AB7";
		s_E349_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AB9";
		s_E350_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ABB";
		s_E351_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ABD";
		s_E352_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ABF";
		s_E353_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AC1";
		s_E354_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AC3";
		s_E355_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AC5";
		s_E356_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AC7";
		s_E357_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AC9";
		s_E358_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ACB";
		s_E359_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ACD";
		s_E360_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ACF";
		s_E361_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AD1";
		s_E362_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AD3";
		s_E363_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AD5";
		s_E364_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AD7";
		s_E365_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AD9";
		s_E366_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ADB";
		s_E367_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ADD";
		s_E368_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ADF";
		s_E369_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AE1";
		s_E370_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AE3";
		s_E371_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AE5";
		s_E372_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AE7";
		s_E373_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AE9";
		s_E374_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AEB";
		s_E375_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AED";
		s_E376_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AEF";
		s_E377_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AF1";
		s_E378_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AF3";
		s_E379_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AF5";
		s_E380_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AF7";
		s_E381_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AF9";
		s_E382_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AFB";
		s_E383_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AFD";
		s_E384_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AFF";
		s_E385_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B01";
		s_E386_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B03";
		s_E387_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B05";
		s_E388_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B07";
		s_E389_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B09";
		s_E390_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B0B";
		s_E391_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B0D";
		s_E392_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B0F";
		s_E393_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B11";
		s_E394_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B13";
		s_E395_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B15";
		s_E396_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B17";
		s_E397_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B19";
		s_E398_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B1B";
		s_E399_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B1D";
		s_E400_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B1F";
		s_E401_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B21";
		s_E402_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B23";
		s_E403_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B25";
		s_E404_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B27";
		s_E405_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B29";
		s_E406_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B2B";
		s_E407_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B2D";
		s_E408_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B2F";
		s_E409_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B31";
		s_E410_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B33";
		s_E411_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B35";
		s_E412_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B37";
		s_E413_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B39";
		s_E414_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B3B";
		s_E415_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B3D";
		s_E416_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B3F";
		s_E417_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B41";
		s_E418_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B43";
		s_E419_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B45";
		s_E420_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B47";
		s_E421_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B49";
		s_E422_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B4B";
		s_E423_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B4D";
		s_E424_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B4F";
		s_E425_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B51";
		s_E426_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B53";
		s_E427_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B55";
		s_E428_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B57";
		s_E429_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B59";
		s_E430_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B5B";
		s_E431_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B5D";
		s_E432_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B5F";
		s_E433_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B61";
		s_E434_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B63";
		s_E435_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B65";
		s_E436_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B67";
		s_E437_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B69";
		s_E438_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B6B";
		s_E439_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B6D";
		s_E440_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B6F";
		s_E441_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B71";
		s_E442_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B73";
		s_E443_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B75";
		s_E444_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B77";
		s_E445_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B79";
		s_E446_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B7B";
		s_E447_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B7D";
		s_E448_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B7F";
		s_E449_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B81";
		s_E450_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B83";
		s_E451_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B85";
		s_E452_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B87";
		s_E453_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B89";
		s_E454_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B8B";
		s_E455_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B8D";
		s_E456_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B8F";
		s_E457_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B91";
		s_E458_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B93";
		s_E459_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B95";
		s_E460_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B97";
		s_E461_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B99";
		s_E462_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B9B";
		s_E463_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B9D";
		s_E464_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B9F";
		s_E465_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BA1";
		s_E466_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BA3";
		s_E467_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BA5";
		s_E468_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BA7";
		s_E469_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BA9";
		s_E470_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BAB";
		s_E471_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BAD";
		s_E472_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BAF";
		s_E473_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BB1";
		s_E474_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BB3";
		s_E475_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BB5";
		s_E476_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BB7";
		s_E477_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BB9";
		s_E478_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BBB";
		s_E479_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BBD";
		s_E480_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BBF";
		s_E481_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BC1";
		s_E482_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BC3";
		s_E483_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BC5";
		s_E484_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BC7";
		s_E485_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BC9";
		s_E486_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BCB";
		s_E487_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BCD";
		s_E488_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BCF";
		s_E489_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BD1";
		s_E490_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BD3";
		s_E491_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BD5";
		s_E492_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BD7";
		s_E493_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BD9";
		s_E494_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BDB";
		s_E495_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BDD";
		s_E496_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BDF";
		s_E497_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BE1";
		s_E498_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BE3";
		s_E499_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BE5";
		s_E500_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BE7";
		s_E501_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BE9";
		s_E502_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BEB";
		s_E503_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BED";
		s_E504_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BEF";
		s_E505_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BF1";
		s_E506_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BF3";
		s_E507_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BF5";
		s_E508_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BF7";
		s_E509_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BF9";
		s_E510_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BFB";
		s_E511_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BFD";
		s_E512_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BFF";
		s_E513_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C01";
		s_E514_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C03";
		s_E515_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C05";
		s_E516_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C07";
		s_E517_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C09";
		s_E518_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C0B";
		s_E519_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C0D";
		s_E520_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C0F";
		s_E521_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C11";
		s_E522_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C13";
		s_E523_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C15";
		s_E524_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C17";
		s_E525_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C19";
		s_E526_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C1B";
		s_E527_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C1D";
		s_E528_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C1F";
		s_E529_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C21";
		s_E530_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C23";
		s_E531_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C25";
		s_E532_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C27";
		s_E533_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C29";
		s_E534_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C2B";
		s_E535_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C2D";
		s_E536_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C2F";
		s_E537_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C31";
		s_E538_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C33";
		s_E539_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C35";
		s_E540_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C37";
		s_E541_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C39";
		s_E542_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C3B";
		s_E543_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C3D";
		s_E544_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C3F";
		s_E545_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C41";
		s_E546_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C43";
		s_E547_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C45";
		s_E548_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C47";
		s_E549_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C49";
		s_E550_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C4B";
		s_E551_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C4D";
		s_E552_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C4F";
		s_E553_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C51";
		s_E554_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C53";
		s_E555_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C55";
		s_E556_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C57";
		s_E557_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C59";
		s_E558_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C5B";
		s_E559_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C5D";
		s_E560_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C5F";
		s_E561_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C61";
		s_E562_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C63";
		s_E563_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C65";
		s_E564_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C67";
		s_E565_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C69";
		s_E566_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C6B";
		s_E567_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C6D";
		s_E568_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C6F";
		s_E569_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C71";
		s_E570_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C73";
		s_E571_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C75";
		s_E572_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C77";
		s_E573_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C79";
		s_E574_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C7B";
		s_E575_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C7D";
		s_E576_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C7F";
		s_E577_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C81";
		s_E578_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C83";
		s_E579_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C85";
		s_E580_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C87";
		s_E581_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C89";
		s_E582_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C8B";
		s_E583_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C8D";
		s_E584_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C8F";
		s_E585_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C91";
		s_E586_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C93";
		s_E587_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C95";
		s_E588_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C97";
		s_E589_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C99";
		s_E590_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C9B";
		s_E591_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C9D";
		s_E592_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C9F";
		s_E593_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CA1";
		s_E594_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CA3";
		s_E595_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CA5";
		s_E596_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CA7";
		s_E597_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CA9";
		s_E598_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CAB";
		s_E599_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CAD";
		s_E600_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CAF";
		s_E601_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CB1";
		s_E602_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CB3";
		s_E603_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CB5";
		s_E604_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CB7";
		s_E605_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CB9";
		s_E606_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CBB";
		s_E607_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CBD";
		s_E608_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CBF";
		s_E609_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CC1";
		s_E610_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CC3";
		s_E611_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CC5";
		s_E612_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CC7";
		s_E613_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CC9";
		s_E614_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CCB";
		s_E615_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CCD";
		s_E616_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CCF";
		s_E617_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CD1";
		s_E618_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CD3";
		s_E619_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CD5";
		s_E620_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CD7";
		s_E621_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CD9";
		s_E622_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CDB";
		s_E623_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CDD";
		s_E624_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CDF";
		s_E625_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CE1";
		s_E626_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CE3";
		s_E627_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CE5";
		s_E628_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CE7";
		s_E629_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CE9";
		s_E630_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CEB";
		s_E631_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CED";
		s_E632_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CEF";
		s_E633_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CF1";
		s_E634_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CF3";
		s_E635_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CF5";
		s_E636_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CF7";
		s_E637_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CF9";
		s_E638_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CFB";
		s_E639_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CFD";
		s_E640_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CFF";
		s_E641_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D01";
		s_E642_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D03";
		s_E643_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D05";
		s_E644_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D07";
		s_E645_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D09";
		s_E646_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D0B";
		s_E647_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D0D";
		s_E648_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D0F";
		s_E649_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D11";
		s_E650_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D13";
		s_E651_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D15";
		s_E652_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D17";
		s_E653_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D19";
		s_E654_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D1B";
		s_E655_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D1D";
		s_E656_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D1F";
		s_E657_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D21";
		s_E658_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D23";
		s_E659_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D25";
		s_E660_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D27";
		s_E661_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D29";
		s_E662_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D2B";
		s_E663_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D2D";
		s_E664_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D2F";
		s_E665_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D31";
		s_E666_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D33";
		s_E667_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D35";
		s_E668_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D37";
		s_E669_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D39";
		s_E670_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D3B";
		s_E671_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D3D";
		s_E672_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D3F";
		s_E673_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D41";
		s_E674_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D43";
		s_E675_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D45";
		s_E676_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D47";
		s_E677_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D49";
		s_E678_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D4B";
		s_E679_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D4D";
		s_E680_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D4F";
		s_E681_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D51";
		s_E682_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D53";
		s_E683_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D55";
		s_E684_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D57";
		s_E685_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D59";
		s_E686_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D5B";
		s_E687_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D5D";
		s_E688_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D5F";
		s_E689_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D61";
		s_E690_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D63";
		s_E691_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D65";
		s_E692_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D67";
		s_E693_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D69";
		s_E694_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D6B";
		s_E695_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D6D";
		s_E696_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D6F";
		s_E697_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D71";
		s_E698_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D73";
		s_E699_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D75";
		s_E700_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D77";
		s_E701_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D79";
		s_E702_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D7B";
		s_E703_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D7D";
		s_E704_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D7F";
		s_E705_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D81";
		s_E706_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D83";
		s_E707_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D85";
		s_E708_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D87";
		s_E709_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D89";
		s_E710_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D8B";
		s_E711_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D8D";
		s_E712_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D8F";
		s_E713_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D91";
		s_E714_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D93";
		s_E715_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D95";
		s_E716_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D97";
		s_E717_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D99";
		s_E718_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D9B";
		s_E719_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D9D";
		s_E720_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D9F";
		s_E721_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DA1";
		s_E722_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DA3";
		s_E723_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DA5";
		s_E724_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DA7";
		s_E725_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DA9";
		s_E726_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DAB";
		s_E727_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DAD";
		s_E728_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DAF";
		s_E729_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DB1";
		s_E730_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DB3";
		s_E731_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DB5";
		s_E732_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DB7";
		s_E733_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DB9";
		s_E734_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DBB";
		s_E735_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DBD";
		s_E736_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DBF";
		s_E737_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DC1";
		s_E738_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DC3";
		s_E739_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DC5";
		s_E740_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DC7";
		s_E741_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DC9";
		s_E742_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DCB";
		s_E743_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DCD";
		s_E744_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DCF";
		s_E745_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DD1";
		s_E746_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DD3";
		s_E747_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DD5";
		s_E748_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DD7";
		s_E749_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DD9";
		s_E750_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DDB";
		s_E751_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DDD";
		s_E752_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DDF";
		s_E753_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DE1";
		s_E754_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DE3";
		s_E755_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DE5";
		s_E756_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DE7";
		s_E757_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DE9";
		s_E758_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DEB";
		s_E759_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DED";
		s_E760_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DEF";
		s_E761_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DF1";
		s_E762_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DF3";
		s_E763_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DF5";
		s_E764_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DF7";
		s_E765_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DF9";
		s_E766_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DFB";
		s_E767_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DFD";
		s_E768_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DFF";
		s_E769_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E01";
		s_E770_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E03";
		s_E771_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E05";
		s_E772_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E07";
		s_E773_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E09";
		s_E774_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E0B";
		s_E775_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E0D";
		s_E776_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E0F";
		s_E777_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E11";
		s_E778_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E13";
		s_E779_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E15";
		s_E780_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E17";
		s_E781_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E19";
		s_E782_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E1B";
		s_E783_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E1D";
		s_E784_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E1F";
		s_E785_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E21";
		s_E786_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E23";
		s_E787_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E25";
		s_E788_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E27";
		s_E789_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E29";
		s_E790_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E2B";
		s_E791_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E2D";
		s_E792_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E2F";
		s_E793_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E31";
		s_E794_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E33";
		s_E795_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E35";
		s_E796_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E37";
		s_E797_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E39";
		s_E798_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E3B";
		s_E799_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E3D";
		s_E800_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E3F";
		s_E801_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E41";
		s_E802_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E43";
		s_E803_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E45";
		s_E804_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E47";
		s_E805_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E49";
		s_E806_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E4B";
		s_E807_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E4D";
		s_E808_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E4F";
		s_E809_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E51";
		s_E810_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E53";
		s_E811_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E55";
		s_E812_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E57";
		s_E813_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E59";
		s_E814_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E5B";
		s_E815_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E5D";
		s_E816_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E5F";
		s_E817_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E61";
		s_E818_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E63";
		s_E819_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E65";
		s_E820_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E67";
		s_E821_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E69";
		s_E822_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E6B";
		s_E823_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E6D";
		s_E824_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E6F";
		s_E825_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E71";
		s_E826_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E73";
		s_E827_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E75";
		s_E828_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E77";
		s_E829_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E79";
		s_E830_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E7B";
		s_E831_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E7D";
		s_E832_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E7F";
		s_E833_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E81";
		s_E834_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E83";
		s_E835_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E85";
		s_E836_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E87";
		s_E837_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E89";
		s_E838_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E8B";
		s_E839_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E8D";
		s_E840_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E8F";
		s_E841_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E91";
		s_E842_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E93";
		s_E843_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E95";
		s_E844_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E97";
		s_E845_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E99";
		s_E846_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E9B";
		s_E847_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E9D";
		s_E848_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E9F";
		s_E849_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EA1";
		s_E850_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EA3";
		s_E851_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EA5";
		s_E852_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EA7";
		s_E853_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EA9";
		s_E854_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EAB";
		s_E855_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EAD";
		s_E856_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EAF";
		s_E857_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EB1";
		s_E858_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EB3";
		s_E859_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EB5";
		s_E860_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EB7";
		s_E861_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EB9";
		s_E862_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EBB";
		s_E863_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EBD";
		s_E864_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EBF";
		s_E865_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EC1";
		s_E866_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EC3";
		s_E867_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EC5";
		s_E868_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EC7";
		s_E869_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EC9";
		s_E870_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ECB";
		s_E871_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ECD";
		s_E872_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ECF";
		s_E873_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ED1";
		s_E874_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ED3";
		s_E875_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ED5";
		s_E876_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ED7";
		s_E877_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ED9";
		s_E878_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EDB";
		s_E879_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EDD";
		s_E880_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EDF";
		s_E881_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EE1";
		s_E882_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EE3";
		s_E883_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EE5";
		s_E884_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EE7";
		s_E885_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EE9";
		s_E886_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EEB";
		s_E887_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EED";
		s_E888_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EEF";
		s_E889_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EF1";
		s_E890_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EF3";
		s_E891_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EF5";
		s_E892_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EF7";
		s_E893_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EF9";
		s_E894_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EFB";
		s_E895_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EFD";
		s_E896_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EFF";
		s_E897_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F01";
		s_E898_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F03";
		s_E899_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F05";
		s_E900_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F07";
		s_E901_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F09";
		s_E902_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F0B";
		s_E903_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F0D";
		s_E904_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F0F";
		s_E905_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F11";
		s_E906_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F13";
		s_E907_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F15";
		s_E908_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F17";
		s_E909_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F19";
		s_E910_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F1B";
		s_E911_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F1D";
		s_E912_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F1F";
		s_E913_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F21";
		s_E914_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F23";
		s_E915_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F25";
		s_E916_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F27";
		s_E917_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F29";
		s_E918_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F2B";
		s_E919_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F2D";
		s_E920_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F2F";
		s_E921_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F31";
		s_E922_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F33";
		s_E923_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F35";
		s_E924_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F37";
		s_E925_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F39";
		s_E926_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F3B";
		s_E927_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F3D";
		s_E928_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F3F";
		s_E929_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F41";
		s_E930_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F43";
		s_E931_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F45";
		s_E932_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F47";
		s_E933_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F49";
		s_E934_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F4B";
		s_E935_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F4D";
		s_E936_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F4F";
		s_E937_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F51";
		s_E938_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F53";
		s_E939_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F55";
		s_E940_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F57";
		s_E941_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F59";
		s_E942_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F5B";
		s_E943_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F5D";
		s_E944_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F5F";
		s_E945_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F61";
		s_E946_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F63";
		s_E947_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F65";
		s_E948_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F67";
		s_E949_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F69";
		s_E950_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F6B";
		s_E951_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F6D";
		s_E952_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F6F";
		s_E953_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F71";
		s_E954_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F73";
		s_E955_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F75";
		s_E956_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F77";
		s_E957_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F79";
		s_E958_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F7B";
		s_E959_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F7D";
		s_E960_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F7F";
		s_E961_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F81";
		s_E962_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F83";
		s_E963_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F85";
		s_E964_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F87";
		s_E965_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F89";
		s_E966_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F8B";
		s_E967_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F8D";
		s_E968_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F8F";
		s_E969_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F91";
		s_E970_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F93";
		s_E971_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F95";
		s_E972_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F97";
		s_E973_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F99";
		s_E974_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F9B";
		s_E975_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F9D";
		s_E976_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F9F";
		s_E977_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FA1";
		s_E978_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FA3";
		s_E979_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FA5";
		s_E980_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FA7";
		s_E981_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FA9";
		s_E982_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FAB";
		s_E983_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FAD";
		s_E984_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FAF";
		s_E985_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FB1";
		s_E986_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FB3";
		s_E987_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FB5";
		s_E988_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FB7";
		s_E989_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FB9";
		s_E990_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FBB";
		s_E991_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FBD";
		s_E992_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FBF";
		s_E993_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FC1";
		s_E994_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FC3";
		s_E995_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FC5";
		s_E996_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FC7";
		s_E997_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FC9";
		s_E998_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FCB";
		s_E999_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FCD";
		s_E1000_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FCF";
		s_E1001_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FD1";
		s_E1002_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FD3";
		s_E1003_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FD5";
		s_E1004_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FD7";
		s_E1005_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FD9";
		s_E1006_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FDB";
		s_E1007_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FDD";
		s_E1008_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FDF";
		s_E1009_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FE1";
		s_E1010_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FE3";
		s_E1011_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FE5";
		s_E1012_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FE7";
		s_E1013_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FE9";
		s_E1014_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FEB";
		s_E1015_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FED";
		s_E1016_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FEF";
		s_E1017_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FF1";
		s_E1018_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FF3";
		s_E1019_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FF5";
		s_E1020_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FF7";
		s_E1021_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FF9";
		s_E1022_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FFB";
		s_E1023_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FFD";
		s_E1024_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FFF";

		s_E2_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"801";
		s_E3_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"803";
		s_E4_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"805";
		s_E5_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"807";
		s_E6_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"809";
		s_E7_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"80B";
		s_E8_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"80D";
		s_E9_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"80F";
		s_E10_C1_L_Pos       	  :std_logic_vector(11 downto 0) := x"811";
		s_E11_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"813";
		s_E12_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"815";
		s_E13_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"817";
		s_E14_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"819";
		s_E15_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"81B";
		s_E16_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"81D";
		s_E17_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"81F";
		s_E18_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"821";
		s_E19_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"823";
		s_E20_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"825";
		s_E21_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"827";
		s_E22_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"829";
		s_E23_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"82B";
		s_E24_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"82D";
		s_E25_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"82F";
		s_E26_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"831";
		s_E27_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"833";
		s_E28_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"835";
		s_E29_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"837";
		s_E30_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"839";
		s_E31_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"83B";
		s_E32_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"83D";
		s_E33_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"83F";
		s_E34_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"841";
		s_E35_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"843";
		s_E36_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"845";
		s_E37_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"847";
		s_E38_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"849";
		s_E39_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"84B";
		s_E40_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"84D";
		s_E41_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"84F";
		s_E42_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"851";
		s_E43_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"853";
		s_E44_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"855";
		s_E45_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"857";
		s_E46_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"859";
		s_E47_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"85B";
		s_E48_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"85D";
		s_E49_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"85F";
		s_E50_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"861";
		s_E51_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"863";
		s_E52_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"865";
		s_E53_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"867";
		s_E54_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"869";
		s_E55_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"86B";
		s_E56_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"86D";
		s_E57_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"86F";
		s_E58_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"871";
		s_E59_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"873";
		s_E60_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"875";
		s_E61_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"877";
		s_E62_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"879";
		s_E63_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"87B";
		s_E64_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"87D";
		s_E65_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"87F";
		s_E66_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"881";
		s_E67_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"883";
		s_E68_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"885";
		s_E69_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"887";
		s_E70_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"889";
		s_E71_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"88B";
		s_E72_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"88D";
		s_E73_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"88F";
		s_E74_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"891";
		s_E75_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"893";
		s_E76_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"895";
		s_E77_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"897";
		s_E78_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"899";
		s_E79_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"89B";
		s_E80_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"89D";
		s_E81_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"89F";
		s_E82_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8A1";
		s_E83_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8A3";
		s_E84_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8A5";
		s_E85_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8A7";
		s_E86_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8A9";
		s_E87_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8AB";
		s_E88_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8AD";
		s_E89_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8AF";
		s_E90_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8B1";
		s_E91_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8B3";
		s_E92_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8B5";
		s_E93_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8B7";
		s_E94_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8B9";
		s_E95_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8BB";
		s_E96_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8BD";
		s_E97_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8BF";
		s_E98_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8C1";
		s_E99_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8C3";
		s_E100_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8C5";
		s_E101_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8C7";
		s_E102_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8C9";
		s_E103_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8CB";
		s_E104_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8CD";
		s_E105_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8CF";
		s_E106_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8D1";
		s_E107_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8D3";
		s_E108_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8D5";
		s_E109_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8D7";
		s_E110_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8D9";
		s_E111_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8DB";
		s_E112_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8DD";
		s_E113_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8DF";
		s_E114_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8E1";
		s_E115_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8E3";
		s_E116_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8E5";
		s_E117_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8E7";
		s_E118_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8E9";
		s_E119_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8EB";
		s_E120_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8ED";
		s_E121_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8EF";
		s_E122_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8F1";
		s_E123_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8F3";
		s_E124_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8F5";
		s_E125_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8F7";
		s_E126_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8F9";
		s_E127_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8FB";
		s_E128_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8FD";
		s_E129_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8FF";
		s_E130_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"901";
		s_E131_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"903";
		s_E132_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"905";
		s_E133_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"907";
		s_E134_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"909";
		s_E135_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"90B";
		s_E136_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"90D";
		s_E137_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"90F";
		s_E138_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"911";
		s_E139_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"913";
		s_E140_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"915";
		s_E141_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"917";
		s_E142_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"919";
		s_E143_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"91B";
		s_E144_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"91D";
		s_E145_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"91F";
		s_E146_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"921";
		s_E147_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"923";
		s_E148_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"925";
		s_E149_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"927";
		s_E150_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"929";
		s_E151_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"92B";
		s_E152_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"92D";
		s_E153_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"92F";
		s_E154_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"931";
		s_E155_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"933";
		s_E156_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"935";
		s_E157_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"937";
		s_E158_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"939";
		s_E159_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"93B";
		s_E160_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"93D";
		s_E161_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"93F";
		s_E162_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"941";
		s_E163_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"943";
		s_E164_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"945";
		s_E165_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"947";
		s_E166_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"949";
		s_E167_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"94B";
		s_E168_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"94D";
		s_E169_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"94F";
		s_E170_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"951";
		s_E171_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"953";
		s_E172_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"955";
		s_E173_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"957";
		s_E174_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"959";
		s_E175_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"95B";
		s_E176_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"95D";
		s_E177_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"95F";
		s_E178_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"961";
		s_E179_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"963";
		s_E180_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"965";
		s_E181_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"967";
		s_E182_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"969";
		s_E183_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"96B";
		s_E184_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"96D";
		s_E185_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"96F";
		s_E186_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"971";
		s_E187_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"973";
		s_E188_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"975";
		s_E189_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"977";
		s_E190_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"979";
		s_E191_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"97B";
		s_E192_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"97D";
		s_E193_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"97F";
		s_E194_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"981";
		s_E195_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"983";
		s_E196_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"985";
		s_E197_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"987";
		s_E198_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"989";
		s_E199_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"98B";
		s_E200_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"98D";
		s_E201_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"98F";
		s_E202_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"991";
		s_E203_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"993";
		s_E204_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"995";
		s_E205_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"997";
		s_E206_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"999";
		s_E207_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"99B";
		s_E208_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"99D";
		s_E209_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"99F";
		s_E210_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9A1";
		s_E211_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9A3";
		s_E212_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9A5";
		s_E213_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9A7";
		s_E214_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9A9";
		s_E215_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9AB";
		s_E216_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9AD";
		s_E217_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9AF";
		s_E218_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9B1";
		s_E219_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9B3";
		s_E220_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9B5";
		s_E221_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9B7";
		s_E222_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9B9";
		s_E223_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9BB";
		s_E224_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9BD";
		s_E225_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9BF";
		s_E226_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9C1";
		s_E227_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9C3";
		s_E228_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9C5";
		s_E229_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9C7";
		s_E230_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9C9";
		s_E231_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9CB";
		s_E232_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9CD";
		s_E233_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9CF";
		s_E234_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9D1";
		s_E235_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9D3";
		s_E236_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9D5";
		s_E237_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9D7";
		s_E238_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9D9";
		s_E239_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9DB";
		s_E240_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9DD";
		s_E241_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9DF";
		s_E242_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9E1";
		s_E243_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9E3";
		s_E244_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9E5";
		s_E245_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9E7";
		s_E246_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9E9";
		s_E247_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9EB";
		s_E248_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9ED";
		s_E249_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9EF";
		s_E250_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9F1";
		s_E251_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9F3";
		s_E252_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9F5";
		s_E253_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9F7";
		s_E254_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9F9";
		s_E255_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9FB";
		s_E256_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9FD";
		s_E257_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9FF";
		s_E258_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A01";
		s_E259_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A03";
		s_E260_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A05";
		s_E261_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A07";
		s_E262_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A09";
		s_E263_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A0B";
		s_E264_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A0D";
		s_E265_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A0F";
		s_E266_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A11";
		s_E267_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A13";
		s_E268_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A15";
		s_E269_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A17";
		s_E270_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A19";
		s_E271_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A1B";
		s_E272_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A1D";
		s_E273_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A1F";
		s_E274_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A21";
		s_E275_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A23";
		s_E276_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A25";
		s_E277_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A27";
		s_E278_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A29";
		s_E279_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A2B";
		s_E280_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A2D";
		s_E281_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A2F";
		s_E282_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A31";
		s_E283_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A33";
		s_E284_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A35";
		s_E285_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A37";
		s_E286_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A39";
		s_E287_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A3B";
		s_E288_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A3D";
		s_E289_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A3F";
		s_E290_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A41";
		s_E291_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A43";
		s_E292_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A45";
		s_E293_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A47";
		s_E294_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A49";
		s_E295_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A4B";
		s_E296_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A4D";
		s_E297_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A4F";
		s_E298_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A51";
		s_E299_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A53";
		s_E300_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A55";
		s_E301_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A57";
		s_E302_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A59";
		s_E303_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A5B";
		s_E304_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A5D";
		s_E305_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A5F";
		s_E306_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A61";
		s_E307_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A63";
		s_E308_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A65";
		s_E309_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A67";
		s_E310_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A69";
		s_E311_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A6B";
		s_E312_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A6D";
		s_E313_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A6F";
		s_E314_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A71";
		s_E315_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A73";
		s_E316_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A75";
		s_E317_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A77";
		s_E318_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A79";
		s_E319_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A7B";
		s_E320_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A7D";
		s_E321_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A7F";
		s_E322_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A81";
		s_E323_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A83";
		s_E324_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A85";
		s_E325_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A87";
		s_E326_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A89";
		s_E327_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A8B";
		s_E328_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A8D";
		s_E329_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A8F";
		s_E330_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A91";
		s_E331_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A93";
		s_E332_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A95";
		s_E333_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A97";
		s_E334_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A99";
		s_E335_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A9B";
		s_E336_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A9D";
		s_E337_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A9F";
		s_E338_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AA1";
		s_E339_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AA3";
		s_E340_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AA5";
		s_E341_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AA7";
		s_E342_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AA9";
		s_E343_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AAB";
		s_E344_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AAD";
		s_E345_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AAF";
		s_E346_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AB1";
		s_E347_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AB3";
		s_E348_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AB5";
		s_E349_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AB7";
		s_E350_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AB9";
		s_E351_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ABB";
		s_E352_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ABD";
		s_E353_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ABF";
		s_E354_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AC1";
		s_E355_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AC3";
		s_E356_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AC5";
		s_E357_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AC7";
		s_E358_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AC9";
		s_E359_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ACB";
		s_E360_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ACD";
		s_E361_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ACF";
		s_E362_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AD1";
		s_E363_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AD3";
		s_E364_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AD5";
		s_E365_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AD7";
		s_E366_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AD9";
		s_E367_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ADB";
		s_E368_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ADD";
		s_E369_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ADF";
		s_E370_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AE1";
		s_E371_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AE3";
		s_E372_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AE5";
		s_E373_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AE7";
		s_E374_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AE9";
		s_E375_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AEB";
		s_E376_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AED";
		s_E377_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AEF";
		s_E378_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AF1";
		s_E379_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AF3";
		s_E380_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AF5";
		s_E381_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AF7";
		s_E382_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AF9";
		s_E383_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AFB";
		s_E384_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AFD";
		s_E385_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AFF";
		s_E386_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B01";
		s_E387_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B03";
		s_E388_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B05";
		s_E389_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B07";
		s_E390_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B09";
		s_E391_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B0B";
		s_E392_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B0D";
		s_E393_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B0F";
		s_E394_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B11";
		s_E395_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B13";
		s_E396_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B15";
		s_E397_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B17";
		s_E398_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B19";
		s_E399_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B1B";
		s_E400_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B1D";
		s_E401_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B1F";
		s_E402_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B21";
		s_E403_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B23";
		s_E404_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B25";
		s_E405_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B27";
		s_E406_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B29";
		s_E407_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B2B";
		s_E408_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B2D";
		s_E409_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B2F";
		s_E410_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B31";
		s_E411_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B33";
		s_E412_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B35";
		s_E413_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B37";
		s_E414_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B39";
		s_E415_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B3B";
		s_E416_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B3D";
		s_E417_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B3F";
		s_E418_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B41";
		s_E419_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B43";
		s_E420_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B45";
		s_E421_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B47";
		s_E422_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B49";
		s_E423_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B4B";
		s_E424_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B4D";
		s_E425_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B4F";
		s_E426_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B51";
		s_E427_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B53";
		s_E428_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B55";
		s_E429_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B57";
		s_E430_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B59";
		s_E431_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B5B";
		s_E432_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B5D";
		s_E433_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B5F";
		s_E434_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B61";
		s_E435_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B63";
		s_E436_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B65";
		s_E437_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B67";
		s_E438_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B69";
		s_E439_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B6B";
		s_E440_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B6D";
		s_E441_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B6F";
		s_E442_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B71";
		s_E443_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B73";
		s_E444_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B75";
		s_E445_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B77";
		s_E446_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B79";
		s_E447_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B7B";
		s_E448_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B7D";
		s_E449_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B7F";
		s_E450_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B81";
		s_E451_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B83";
		s_E452_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B85";
		s_E453_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B87";
		s_E454_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B89";
		s_E455_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B8B";
		s_E456_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B8D";
		s_E457_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B8F";
		s_E458_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B91";
		s_E459_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B93";
		s_E460_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B95";
		s_E461_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B97";
		s_E462_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B99";
		s_E463_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B9B";
		s_E464_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B9D";
		s_E465_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B9F";
		s_E466_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BA1";
		s_E467_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BA3";
		s_E468_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BA5";
		s_E469_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BA7";
		s_E470_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BA9";
		s_E471_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BAB";
		s_E472_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BAD";
		s_E473_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BAF";
		s_E474_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BB1";
		s_E475_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BB3";
		s_E476_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BB5";
		s_E477_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BB7";
		s_E478_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BB9";
		s_E479_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BBB";
		s_E480_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BBD";
		s_E481_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BBF";
		s_E482_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BC1";
		s_E483_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BC3";
		s_E484_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BC5";
		s_E485_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BC7";
		s_E486_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BC9";
		s_E487_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BCB";
		s_E488_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BCD";
		s_E489_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BCF";
		s_E490_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BD1";
		s_E491_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BD3";
		s_E492_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BD5";
		s_E493_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BD7";
		s_E494_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BD9";
		s_E495_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BDB";
		s_E496_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BDD";
		s_E497_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BDF";
		s_E498_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BE1";
		s_E499_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BE3";
		s_E500_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BE5";
		s_E501_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BE7";
		s_E502_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BE9";
		s_E503_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BEB";
		s_E504_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BED";
		s_E505_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BEF";
		s_E506_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BF1";
		s_E507_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BF3";
		s_E508_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BF5";
		s_E509_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BF7";
		s_E510_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BF9";
		s_E511_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BFB";
		s_E512_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BFD";
		s_E513_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BFF";
		s_E514_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C01";
		s_E515_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C03";
		s_E516_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C05";
		s_E517_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C07";
		s_E518_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C09";
		s_E519_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C0B";
		s_E520_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C0D";
		s_E521_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C0F";
		s_E522_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C11";
		s_E523_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C13";
		s_E524_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C15";
		s_E525_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C17";
		s_E526_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C19";
		s_E527_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C1B";
		s_E528_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C1D";
		s_E529_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C1F";
		s_E530_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C21";
		s_E531_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C23";
		s_E532_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C25";
		s_E533_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C27";
		s_E534_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C29";
		s_E535_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C2B";
		s_E536_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C2D";
		s_E537_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C2F";
		s_E538_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C31";
		s_E539_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C33";
		s_E540_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C35";
		s_E541_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C37";
		s_E542_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C39";
		s_E543_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C3B";
		s_E544_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C3D";
		s_E545_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C3F";
		s_E546_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C41";
		s_E547_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C43";
		s_E548_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C45";
		s_E549_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C47";
		s_E550_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C49";
		s_E551_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C4B";
		s_E552_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C4D";
		s_E553_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C4F";
		s_E554_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C51";
		s_E555_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C53";
		s_E556_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C55";
		s_E557_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C57";
		s_E558_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C59";
		s_E559_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C5B";
		s_E560_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C5D";
		s_E561_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C5F";
		s_E562_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C61";
		s_E563_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C63";
		s_E564_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C65";
		s_E565_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C67";
		s_E566_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C69";
		s_E567_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C6B";
		s_E568_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C6D";
		s_E569_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C6F";
		s_E570_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C71";
		s_E571_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C73";
		s_E572_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C75";
		s_E573_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C77";
		s_E574_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C79";
		s_E575_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C7B";
		s_E576_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C7D";
		s_E577_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C7F";
		s_E578_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C81";
		s_E579_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C83";
		s_E580_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C85";
		s_E581_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C87";
		s_E582_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C89";
		s_E583_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C8B";
		s_E584_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C8D";
		s_E585_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C8F";
		s_E586_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C91";
		s_E587_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C93";
		s_E588_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C95";
		s_E589_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C97";
		s_E590_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C99";
		s_E591_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C9B";
		s_E592_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C9D";
		s_E593_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C9F";
		s_E594_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CA1";
		s_E595_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CA3";
		s_E596_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CA5";
		s_E597_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CA7";
		s_E598_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CA9";
		s_E599_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CAB";
		s_E600_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CAD";
		s_E601_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CAF";
		s_E602_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CB1";
		s_E603_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CB3";
		s_E604_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CB5";
		s_E605_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CB7";
		s_E606_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CB9";
		s_E607_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CBB";
		s_E608_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CBD";
		s_E609_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CBF";
		s_E610_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CC1";
		s_E611_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CC3";
		s_E612_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CC5";
		s_E613_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CC7";
		s_E614_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CC9";
		s_E615_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CCB";
		s_E616_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CCD";
		s_E617_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CCF";
		s_E618_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CD1";
		s_E619_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CD3";
		s_E620_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CD5";
		s_E621_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CD7";
		s_E622_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CD9";
		s_E623_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CDB";
		s_E624_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CDD";
		s_E625_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CDF";
		s_E626_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CE1";
		s_E627_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CE3";
		s_E628_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CE5";
		s_E629_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CE7";
		s_E630_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CE9";
		s_E631_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CEB";
		s_E632_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CED";
		s_E633_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CEF";
		s_E634_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CF1";
		s_E635_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CF3";
		s_E636_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CF5";
		s_E637_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CF7";
		s_E638_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CF9";
		s_E639_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CFB";
		s_E640_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CFD";
		s_E641_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CFF";
		s_E642_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D01";
		s_E643_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D03";
		s_E644_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D05";
		s_E645_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D07";
		s_E646_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D09";
		s_E647_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D0B";
		s_E648_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D0D";
		s_E649_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D0F";
		s_E650_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D11";
		s_E651_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D13";
		s_E652_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D15";
		s_E653_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D17";
		s_E654_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D19";
		s_E655_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D1B";
		s_E656_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D1D";
		s_E657_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D1F";
		s_E658_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D21";
		s_E659_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D23";
		s_E660_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D25";
		s_E661_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D27";
		s_E662_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D29";
		s_E663_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D2B";
		s_E664_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D2D";
		s_E665_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D2F";
		s_E666_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D31";
		s_E667_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D33";
		s_E668_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D35";
		s_E669_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D37";
		s_E670_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D39";
		s_E671_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D3B";
		s_E672_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D3D";
		s_E673_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D3F";
		s_E674_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D41";
		s_E675_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D43";
		s_E676_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D45";
		s_E677_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D47";
		s_E678_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D49";
		s_E679_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D4B";
		s_E680_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D4D";
		s_E681_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D4F";
		s_E682_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D51";
		s_E683_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D53";
		s_E684_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D55";
		s_E685_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D57";
		s_E686_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D59";
		s_E687_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D5B";
		s_E688_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D5D";
		s_E689_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D5F";
		s_E690_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D61";
		s_E691_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D63";
		s_E692_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D65";
		s_E693_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D67";
		s_E694_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D69";
		s_E695_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D6B";
		s_E696_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D6D";
		s_E697_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D6F";
		s_E698_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D71";
		s_E699_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D73";
		s_E700_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D75";
		s_E701_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D77";
		s_E702_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D79";
		s_E703_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D7B";
		s_E704_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D7D";
		s_E705_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D7F";
		s_E706_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D81";
		s_E707_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D83";
		s_E708_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D85";
		s_E709_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D87";
		s_E710_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D89";
		s_E711_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D8B";
		s_E712_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D8D";
		s_E713_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D8F";
		s_E714_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D91";
		s_E715_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D93";
		s_E716_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D95";
		s_E717_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D97";
		s_E718_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D99";
		s_E719_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D9B";
		s_E720_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D9D";
		s_E721_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D9F";
		s_E722_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DA1";
		s_E723_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DA3";
		s_E724_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DA5";
		s_E725_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DA7";
		s_E726_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DA9";
		s_E727_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DAB";
		s_E728_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DAD";
		s_E729_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DAF";
		s_E730_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DB1";
		s_E731_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DB3";
		s_E732_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DB5";
		s_E733_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DB7";
		s_E734_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DB9";
		s_E735_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DBB";
		s_E736_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DBD";
		s_E737_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DBF";
		s_E738_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DC1";
		s_E739_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DC3";
		s_E740_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DC5";
		s_E741_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DC7";
		s_E742_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DC9";
		s_E743_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DCB";
		s_E744_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DCD";
		s_E745_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DCF";
		s_E746_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DD1";
		s_E747_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DD3";
		s_E748_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DD5";
		s_E749_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DD7";
		s_E750_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DD9";
		s_E751_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DDB";
		s_E752_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DDD";
		s_E753_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DDF";
		s_E754_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DE1";
		s_E755_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DE3";
		s_E756_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DE5";
		s_E757_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DE7";
		s_E758_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DE9";
		s_E759_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DEB";
		s_E760_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DED";
		s_E761_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DEF";
		s_E762_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DF1";
		s_E763_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DF3";
		s_E764_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DF5";
		s_E765_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DF7";
		s_E766_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DF9";
		s_E767_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DFB";
		s_E768_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DFD";
		s_E769_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DFF";
		s_E770_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E01";
		s_E771_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E03";
		s_E772_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E05";
		s_E773_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E07";
		s_E774_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E09";
		s_E775_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E0B";
		s_E776_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E0D";
		s_E777_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E0F";
		s_E778_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E11";
		s_E779_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E13";
		s_E780_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E15";
		s_E781_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E17";
		s_E782_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E19";
		s_E783_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E1B";
		s_E784_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E1D";
		s_E785_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E1F";
		s_E786_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E21";
		s_E787_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E23";
		s_E788_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E25";
		s_E789_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E27";
		s_E790_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E29";
		s_E791_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E2B";
		s_E792_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E2D";
		s_E793_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E2F";
		s_E794_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E31";
		s_E795_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E33";
		s_E796_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E35";
		s_E797_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E37";
		s_E798_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E39";
		s_E799_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E3B";
		s_E800_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E3D";
		s_E801_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E3F";
		s_E802_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E41";
		s_E803_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E43";
		s_E804_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E45";
		s_E805_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E47";
		s_E806_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E49";
		s_E807_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E4B";
		s_E808_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E4D";
		s_E809_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E4F";
		s_E810_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E51";
		s_E811_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E53";
		s_E812_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E55";
		s_E813_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E57";
		s_E814_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E59";
		s_E815_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E5B";
		s_E816_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E5D";
		s_E817_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E5F";
		s_E818_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E61";
		s_E819_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E63";
		s_E820_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E65";
		s_E821_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E67";
		s_E822_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E69";
		s_E823_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E6B";
		s_E824_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E6D";
		s_E825_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E6F";
		s_E826_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E71";
		s_E827_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E73";
		s_E828_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E75";
		s_E829_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E77";
		s_E830_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E79";
		s_E831_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E7B";
		s_E832_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E7D";
		s_E833_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E7F";
		s_E834_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E81";
		s_E835_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E83";
		s_E836_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E85";
		s_E837_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E87";
		s_E838_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E89";
		s_E839_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E8B";
		s_E840_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E8D";
		s_E841_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E8F";
		s_E842_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E91";
		s_E843_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E93";
		s_E844_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E95";
		s_E845_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E97";
		s_E846_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E99";
		s_E847_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E9B";
		s_E848_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E9D";
		s_E849_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E9F";
		s_E850_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EA1";
		s_E851_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EA3";
		s_E852_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EA5";
		s_E853_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EA7";
		s_E854_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EA9";
		s_E855_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EAB";
		s_E856_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EAD";
		s_E857_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EAF";
		s_E858_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EB1";
		s_E859_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EB3";
		s_E860_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EB5";
		s_E861_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EB7";
		s_E862_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EB9";
		s_E863_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EBB";
		s_E864_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EBD";
		s_E865_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EBF";
		s_E866_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EC1";
		s_E867_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EC3";
		s_E868_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EC5";
		s_E869_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EC7";
		s_E870_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EC9";
		s_E871_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ECB";
		s_E872_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ECD";
		s_E873_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ECF";
		s_E874_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ED1";
		s_E875_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ED3";
		s_E876_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ED5";
		s_E877_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ED7";
		s_E878_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ED9";
		s_E879_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EDB";
		s_E880_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EDD";
		s_E881_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EDF";
		s_E882_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EE1";
		s_E883_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EE3";
		s_E884_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EE5";
		s_E885_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EE7";
		s_E886_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EE9";
		s_E887_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EEB";
		s_E888_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EED";
		s_E889_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EEF";
		s_E890_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EF1";
		s_E891_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EF3";
		s_E892_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EF5";
		s_E893_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EF7";
		s_E894_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EF9";
		s_E895_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EFB";
		s_E896_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EFD";
		s_E897_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EFF";
		s_E898_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F01";
		s_E899_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F03";
		s_E900_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F05";
		s_E901_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F07";
		s_E902_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F09";
		s_E903_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F0B";
		s_E904_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F0D";
		s_E905_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F0F";
		s_E906_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F11";
		s_E907_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F13";
		s_E908_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F15";
		s_E909_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F17";
		s_E910_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F19";
		s_E911_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F1B";
		s_E912_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F1D";
		s_E913_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F1F";
		s_E914_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F21";
		s_E915_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F23";
		s_E916_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F25";
		s_E917_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F27";
		s_E918_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F29";
		s_E919_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F2B";
		s_E920_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F2D";
		s_E921_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F2F";
		s_E922_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F31";
		s_E923_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F33";
		s_E924_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F35";
		s_E925_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F37";
		s_E926_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F39";
		s_E927_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F3B";
		s_E928_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F3D";
		s_E929_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F3F";
		s_E930_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F41";
		s_E931_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F43";
		s_E932_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F45";
		s_E933_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F47";
		s_E934_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F49";
		s_E935_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F4B";
		s_E936_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F4D";
		s_E937_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F4F";
		s_E938_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F51";
		s_E939_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F53";
		s_E940_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F55";
		s_E941_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F57";
		s_E942_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F59";
		s_E943_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F5B";
		s_E944_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F5D";
		s_E945_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F5F";
		s_E946_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F61";
		s_E947_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F63";
		s_E948_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F65";
		s_E949_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F67";
		s_E950_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F69";
		s_E951_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F6B";
		s_E952_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F6D";
		s_E953_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F6F";
		s_E954_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F71";
		s_E955_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F73";
		s_E956_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F75";
		s_E957_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F77";
		s_E958_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F79";
		s_E959_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F7B";
		s_E960_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F7D";
		s_E961_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F7F";
		s_E962_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F81";
		s_E963_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F83";
		s_E964_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F85";
		s_E965_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F87";
		s_E966_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F89";
		s_E967_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F8B";
		s_E968_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F8D";
		s_E969_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F8F";
		s_E970_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F91";
		s_E971_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F93";
		s_E972_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F95";
		s_E973_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F97";
		s_E974_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F99";
		s_E975_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F9B";
		s_E976_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F9D";
		s_E977_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F9F";
		s_E978_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FA1";
		s_E979_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FA3";
		s_E980_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FA5";
		s_E981_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FA7";
		s_E982_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FA9";
		s_E983_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FAB";
		s_E984_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FAD";
		s_E985_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FAF";
		s_E986_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FB1";
		s_E987_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FB3";
		s_E988_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FB5";
		s_E989_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FB7";
		s_E990_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FB9";
		s_E991_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FBB";
		s_E992_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FBD";
		s_E993_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FBF";
		s_E994_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FC1";
		s_E995_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FC3";
		s_E996_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FC5";
		s_E997_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FC7";
		s_E998_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FC9";
		s_E999_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FCB";
		s_E1000_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FCD";
		s_E1001_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FCF";
		s_E1002_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FD1";
		s_E1003_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FD3";
		s_E1004_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FD5";
		s_E1005_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FD7";
		s_E1006_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FD9";
		s_E1007_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FDB";
		s_E1008_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FDD";
		s_E1009_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FDF";
		s_E1010_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FE1";
		s_E1011_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FE3";
		s_E1012_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FE5";
		s_E1013_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FE7";
		s_E1014_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FE9";
		s_E1015_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FEB";
		s_E1016_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FED";
		s_E1017_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FEF";
		s_E1018_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FF1";
		s_E1019_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FF3";
		s_E1020_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FF5";
		s_E1021_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FF7";
		s_E1022_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FF9";
		s_E1023_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FFB";
		s_E1024_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FFD"

      );

  --+----------
  -- Port name declarations
  --+----------
  port   (
       CLK100     			   :in  std_logic;
       RST        			   :in  std_logic;
       
       DATA1                   :in  std_logic_vector(WdVecSize_g-5 downto 0);
       DATARDY1                :in  std_logic;
       DATA2                   :in  std_logic_vector(WdVecSize_g-5 downto 0);
       DATARDY2                :in  std_logic;
        
--       THRESHOLD  :in  std_logic_vector(NibbleSize_g-1 downto 0);
       
	   ADD_TIMP_FLAG 		   :out std_logic;
	   ADD_TIMP_FLAG_pos 	   :out std_logic;
	   
	   o_DATA_OUT_C1  		   :out std_logic_vector(11 downto 0);
	   o_DATA_OUT_C2  		   :out std_logic_vector(11 downto 0);
							   
       i_PEAK_THD          	   :in std_logic_vector(11 downto 0);
       i_PEAK_THD_pos          :in std_logic_vector(11 downto 0);

	   o_Energy_Bin_1    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_2    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_3    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_4    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_5    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_6    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_7    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_8    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_9    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_10   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_11   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_12   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_13   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_14   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_15   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_16   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_17   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_18   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_19   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_20   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_21   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_22   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_23   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_24   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_25   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_26   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_27   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_28   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_29   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_30   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_31   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_32   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_33   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_34   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_35   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_36   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_37   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_38   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_39   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_40   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_41   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_42   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_43   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_44   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_45   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_46   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_47   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_48   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_49   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_50   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_51   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_52   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_53   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_54   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_55   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_56   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_57   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_58   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_59   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_60   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_61   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_62   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_63   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_64   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_65   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_66   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_67   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_68   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_69   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_70   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_71   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_72   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_73   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_74   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_75   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_76   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_77   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_78   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_79   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_80   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_81   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_82   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_83   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_84   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_85   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_86   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_87   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_88   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_89   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_90   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_91   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_92   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_93   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_94   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_95   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_96   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_97   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_98   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_99   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_100  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_101  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_102  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_103  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_104  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_105  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_106  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_107  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_108  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_109  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_110  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_111  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_112  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_113  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_114  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_115  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_116  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_117  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_118  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_119  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_120  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_121  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_122  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_123  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_124  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_125  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_126  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_127  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_128  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_129  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_130  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_131  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_132  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_133  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_134  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_135  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_136  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_137  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_138  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_139  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_140  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_141  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_142  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_143  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_144  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_145  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_146  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_147  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_148  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_149  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_150  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_151  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_152  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_153  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_154  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_155  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_156  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_157  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_158  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_159  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_160  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_161  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_162  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_163  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_164  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_165  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_166  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_167  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_168  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_169  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_170  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_171  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_172  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_173  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_174  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_175  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_176  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_177  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_178  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_179  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_180  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_181  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_182  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_183  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_184  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_185  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_186  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_187  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_188  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_189  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_190  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_191  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_192  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_193  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_194  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_195  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_196  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_197  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_198  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_199  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_200  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_201  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_202  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_203  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_204  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_205  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_206  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_207  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_208  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_209  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_210  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_211  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_212  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_213  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_214  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_215  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_216  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_217  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_218  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_219  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_220  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_221  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_222  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_223  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_224  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_225  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_226  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_227  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_228  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_229  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_230  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_231  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_232  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_233  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_234  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_235  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_236  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_237  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_238  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_239  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_240  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_241  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_242  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_243  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_244  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_245  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_246  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_247  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_248  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_249  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_250  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_251  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_252  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_253  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_254  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_255  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_256  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_257  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_258  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_259  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_260  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_261  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_262  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_263  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_264  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_265  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_266  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_267  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_268  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_269  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_270  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_271  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_272  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_273  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_274  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_275  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_276  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_277  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_278  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_279  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_280  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_281  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_282  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_283  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_284  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_285  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_286  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_287  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_288  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_289  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_290  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_291  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_292  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_293  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_294  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_295  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_296  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_297  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_298  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_299  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_300  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_301  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_302  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_303  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_304  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_305  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_306  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_307  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_308  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_309  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_310  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_311  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_312  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_313  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_314  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_315  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_316  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_317  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_318  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_319  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_320  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_321  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_322  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_323  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_324  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_325  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_326  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_327  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_328  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_329  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_330  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_331  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_332  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_333  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_334  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_335  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_336  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_337  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_338  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_339  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_340  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_341  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_342  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_343  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_344  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_345  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_346  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_347  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_348  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_349  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_350  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_351  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_352  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_353  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_354  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_355  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_356  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_357  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_358  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_359  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_360  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_361  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_362  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_363  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_364  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_365  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_366  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_367  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_368  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_369  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_370  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_371  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_372  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_373  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_374  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_375  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_376  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_377  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_378  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_379  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_380  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_381  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_382  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_383  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_384  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_385  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_386  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_387  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_388  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_389  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_390  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_391  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_392  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_393  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_394  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_395  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_396  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_397  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_398  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_399  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_400  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_401  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_402  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_403  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_404  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_405  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_406  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_407  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_408  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_409  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_410  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_411  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_412  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_413  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_414  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_415  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_416  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_417  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_418  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_419  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_420  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_421  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_422  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_423  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_424  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_425  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_426  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_427  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_428  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_429  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_430  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_431  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_432  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_433  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_434  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_435  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_436  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_437  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_438  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_439  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_440  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_441  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_442  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_443  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_444  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_445  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_446  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_447  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_448  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_449  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_450  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_451  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_452  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_453  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_454  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_455  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_456  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_457  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_458  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_459  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_460  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_461  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_462  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_463  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_464  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_465  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_466  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_467  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_468  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_469  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_470  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_471  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_472  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_473  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_474  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_475  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_476  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_477  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_478  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_479  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_480  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_481  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_482  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_483  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_484  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_485  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_486  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_487  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_488  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_489  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_490  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_491  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_492  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_493  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_494  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_495  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_496  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_497  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_498  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_499  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_500  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_501  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_502  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_503  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_504  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_505  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_506  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_507  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_508  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_509  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_510  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_511  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_512  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_513  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_514  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_515  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_516  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_517  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_518  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_519  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_520  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_521  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_522  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_523  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_524  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_525  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_526  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_527  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_528  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_529  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_530  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_531  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_532  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_533  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_534  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_535  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_536  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_537  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_538  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_539  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_540  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_541  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_542  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_543  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_544  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_545  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_546  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_547  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_548  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_549  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_550  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_551  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_552  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_553  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_554  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_555  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_556  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_557  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_558  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_559  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_560  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_561  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_562  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_563  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_564  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_565  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_566  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_567  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_568  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_569  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_570  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_571  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_572  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_573  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_574  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_575  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_576  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_577  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_578  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_579  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_580  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_581  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_582  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_583  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_584  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_585  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_586  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_587  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_588  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_589  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_590  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_591  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_592  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_593  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_594  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_595  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_596  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_597  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_598  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_599  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_600  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_601  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_602  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_603  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_604  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_605  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_606  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_607  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_608  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_609  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_610  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_611  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_612  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_613  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_614  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_615  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_616  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_617  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_618  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_619  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_620  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_621  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_622  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_623  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_624  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_625  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_626  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_627  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_628  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_629  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_630  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_631  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_632  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_633  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_634  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_635  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_636  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_637  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_638  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_639  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_640  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_641  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_642  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_643  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_644  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_645  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_646  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_647  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_648  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_649  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_650  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_651  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_652  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_653  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_654  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_655  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_656  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_657  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_658  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_659  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_660  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_661  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_662  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_663  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_664  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_665  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_666  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_667  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_668  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_669  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_670  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_671  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_672  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_673  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_674  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_675  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_676  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_677  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_678  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_679  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_680  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_681  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_682  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_683  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_684  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_685  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_686  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_687  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_688  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_689  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_690  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_691  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_692  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_693  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_694  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_695  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_696  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_697  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_698  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_699  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_700  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_701  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_702  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_703  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_704  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_705  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_706  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_707  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_708  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_709  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_710  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_711  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_712  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_713  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_714  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_715  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_716  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_717  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_718  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_719  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_720  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_721  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_722  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_723  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_724  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_725  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_726  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_727  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_728  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_729  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_730  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_731  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_732  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_733  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_734  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_735  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_736  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_737  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_738  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_739  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_740  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_741  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_742  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_743  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_744  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_745  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_746  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_747  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_748  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_749  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_750  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_751  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_752  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_753  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_754  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_755  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_756  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_757  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_758  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_759  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_760  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_761  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_762  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_763  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_764  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_765  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_766  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_767  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_768  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_769  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_770  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_771  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_772  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_773  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_774  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_775  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_776  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_777  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_778  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_779  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_780  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_781  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_782  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_783  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_784  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_785  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_786  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_787  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_788  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_789  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_790  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_791  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_792  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_793  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_794  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_795  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_796  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_797  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_798  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_799  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_800  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_801  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_802  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_803  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_804  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_805  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_806  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_807  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_808  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_809  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_810  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_811  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_812  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_813  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_814  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_815  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_816  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_817  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_818  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_819  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_820  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_821  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_822  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_823  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_824  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_825  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_826  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_827  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_828  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_829  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_830  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_831  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_832  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_833  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_834  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_835  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_836  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_837  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_838  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_839  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_840  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_841  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_842  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_843  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_844  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_845  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_846  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_847  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_848  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_849  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_850  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_851  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_852  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_853  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_854  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_855  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_856  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_857  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_858  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_859  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_860  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_861  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_862  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_863  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_864  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_865  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_866  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_867  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_868  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_869  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_870  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_871  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_872  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_873  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_874  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_875  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_876  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_877  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_878  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_879  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_880  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_881  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_882  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_883  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_884  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_885  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_886  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_887  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_888  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_889  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_890  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_891  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_892  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_893  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_894  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_895  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_896  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_897  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_898  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_899  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_900  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_901  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_902  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_903  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_904  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_905  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_906  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_907  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_908  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_909  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_910  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_911  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_912  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_913  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_914  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_915  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_916  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_917  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_918  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_919  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_920  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_921  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_922  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_923  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_924  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_925  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_926  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_927  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_928  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_929  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_930  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_931  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_932  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_933  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_934  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_935  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_936  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_937  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_938  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_939  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_940  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_941  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_942  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_943  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_944  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_945  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_946  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_947  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_948  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_949  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_950  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_951  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_952  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_953  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_954  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_955  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_956  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_957  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_958  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_959  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_960  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_961  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_962  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_963  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_964  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_965  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_966  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_967  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_968  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_969  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_970  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_971  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_972  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_973  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_974  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_975  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_976  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_977  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_978  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_979  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_980  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_981  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_982  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_983  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_984  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_985  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_986  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_987  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_988  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_989  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_990  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_991  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_992  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_993  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_994  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_995  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_996  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_997  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_998  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_999  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1000 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1001 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1002 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1003 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1004 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1005 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1006 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1007 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1008 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1009 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1010 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1011 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1012 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1013 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1014 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1015 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1016 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1017 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1018 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1019 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1020 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1021 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1022 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1023 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1024 :out std_logic_vector(11 downto 0);
	   
	   o_Energy_Bin_Pos_1    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_2    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_3    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_4    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_5    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_6    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_7    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_8    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_9    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_10   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_11   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_12   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_13   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_14   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_15   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_16   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_17   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_18   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_19   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_20   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_21   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_22   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_23   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_24   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_25   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_26   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_27   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_28   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_29   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_30   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_31   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_32   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_33   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_34   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_35   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_36   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_37   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_38   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_39   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_40   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_41   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_42   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_43   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_44   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_45   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_46   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_47   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_48   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_49   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_50   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_51   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_52   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_53   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_54   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_55   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_56   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_57   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_58   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_59   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_60   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_61   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_62   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_63   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_64   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_65   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_66   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_67   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_68   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_69   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_70   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_71   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_72   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_73   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_74   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_75   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_76   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_77   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_78   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_79   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_80   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_81   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_82   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_83   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_84   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_85   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_86   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_87   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_88   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_89   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_90   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_91   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_92   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_93   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_94   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_95   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_96   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_97   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_98   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_99   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_100  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_101  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_102  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_103  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_104  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_105  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_106  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_107  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_108  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_109  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_110  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_111  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_112  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_113  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_114  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_115  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_116  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_117  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_118  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_119  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_120  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_121  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_122  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_123  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_124  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_125  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_126  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_127  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_128  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_129  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_130  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_131  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_132  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_133  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_134  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_135  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_136  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_137  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_138  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_139  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_140  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_141  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_142  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_143  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_144  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_145  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_146  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_147  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_148  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_149  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_150  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_151  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_152  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_153  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_154  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_155  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_156  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_157  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_158  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_159  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_160  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_161  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_162  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_163  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_164  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_165  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_166  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_167  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_168  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_169  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_170  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_171  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_172  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_173  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_174  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_175  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_176  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_177  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_178  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_179  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_180  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_181  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_182  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_183  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_184  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_185  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_186  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_187  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_188  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_189  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_190  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_191  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_192  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_193  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_194  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_195  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_196  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_197  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_198  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_199  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_200  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_201  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_202  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_203  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_204  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_205  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_206  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_207  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_208  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_209  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_210  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_211  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_212  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_213  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_214  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_215  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_216  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_217  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_218  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_219  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_220  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_221  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_222  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_223  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_224  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_225  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_226  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_227  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_228  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_229  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_230  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_231  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_232  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_233  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_234  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_235  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_236  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_237  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_238  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_239  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_240  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_241  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_242  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_243  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_244  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_245  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_246  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_247  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_248  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_249  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_250  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_251  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_252  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_253  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_254  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_255  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_256  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_257  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_258  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_259  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_260  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_261  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_262  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_263  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_264  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_265  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_266  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_267  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_268  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_269  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_270  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_271  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_272  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_273  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_274  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_275  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_276  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_277  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_278  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_279  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_280  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_281  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_282  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_283  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_284  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_285  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_286  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_287  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_288  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_289  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_290  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_291  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_292  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_293  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_294  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_295  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_296  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_297  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_298  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_299  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_300  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_301  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_302  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_303  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_304  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_305  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_306  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_307  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_308  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_309  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_310  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_311  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_312  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_313  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_314  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_315  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_316  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_317  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_318  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_319  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_320  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_321  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_322  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_323  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_324  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_325  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_326  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_327  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_328  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_329  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_330  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_331  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_332  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_333  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_334  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_335  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_336  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_337  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_338  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_339  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_340  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_341  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_342  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_343  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_344  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_345  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_346  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_347  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_348  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_349  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_350  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_351  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_352  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_353  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_354  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_355  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_356  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_357  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_358  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_359  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_360  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_361  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_362  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_363  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_364  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_365  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_366  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_367  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_368  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_369  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_370  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_371  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_372  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_373  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_374  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_375  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_376  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_377  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_378  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_379  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_380  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_381  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_382  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_383  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_384  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_385  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_386  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_387  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_388  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_389  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_390  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_391  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_392  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_393  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_394  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_395  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_396  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_397  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_398  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_399  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_400  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_401  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_402  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_403  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_404  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_405  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_406  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_407  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_408  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_409  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_410  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_411  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_412  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_413  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_414  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_415  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_416  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_417  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_418  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_419  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_420  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_421  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_422  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_423  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_424  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_425  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_426  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_427  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_428  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_429  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_430  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_431  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_432  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_433  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_434  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_435  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_436  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_437  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_438  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_439  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_440  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_441  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_442  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_443  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_444  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_445  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_446  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_447  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_448  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_449  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_450  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_451  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_452  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_453  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_454  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_455  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_456  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_457  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_458  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_459  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_460  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_461  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_462  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_463  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_464  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_465  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_466  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_467  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_468  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_469  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_470  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_471  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_472  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_473  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_474  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_475  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_476  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_477  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_478  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_479  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_480  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_481  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_482  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_483  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_484  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_485  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_486  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_487  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_488  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_489  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_490  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_491  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_492  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_493  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_494  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_495  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_496  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_497  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_498  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_499  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_500  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_501  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_502  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_503  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_504  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_505  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_506  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_507  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_508  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_509  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_510  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_511  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_512  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_513  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_514  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_515  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_516  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_517  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_518  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_519  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_520  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_521  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_522  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_523  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_524  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_525  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_526  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_527  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_528  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_529  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_530  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_531  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_532  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_533  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_534  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_535  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_536  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_537  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_538  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_539  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_540  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_541  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_542  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_543  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_544  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_545  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_546  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_547  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_548  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_549  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_550  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_551  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_552  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_553  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_554  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_555  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_556  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_557  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_558  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_559  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_560  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_561  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_562  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_563  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_564  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_565  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_566  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_567  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_568  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_569  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_570  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_571  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_572  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_573  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_574  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_575  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_576  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_577  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_578  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_579  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_580  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_581  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_582  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_583  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_584  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_585  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_586  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_587  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_588  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_589  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_590  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_591  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_592  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_593  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_594  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_595  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_596  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_597  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_598  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_599  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_600  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_601  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_602  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_603  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_604  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_605  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_606  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_607  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_608  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_609  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_610  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_611  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_612  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_613  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_614  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_615  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_616  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_617  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_618  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_619  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_620  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_621  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_622  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_623  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_624  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_625  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_626  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_627  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_628  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_629  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_630  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_631  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_632  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_633  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_634  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_635  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_636  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_637  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_638  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_639  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_640  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_641  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_642  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_643  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_644  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_645  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_646  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_647  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_648  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_649  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_650  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_651  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_652  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_653  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_654  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_655  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_656  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_657  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_658  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_659  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_660  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_661  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_662  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_663  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_664  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_665  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_666  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_667  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_668  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_669  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_670  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_671  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_672  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_673  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_674  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_675  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_676  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_677  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_678  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_679  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_680  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_681  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_682  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_683  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_684  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_685  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_686  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_687  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_688  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_689  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_690  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_691  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_692  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_693  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_694  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_695  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_696  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_697  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_698  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_699  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_700  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_701  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_702  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_703  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_704  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_705  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_706  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_707  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_708  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_709  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_710  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_711  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_712  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_713  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_714  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_715  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_716  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_717  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_718  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_719  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_720  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_721  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_722  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_723  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_724  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_725  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_726  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_727  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_728  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_729  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_730  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_731  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_732  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_733  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_734  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_735  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_736  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_737  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_738  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_739  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_740  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_741  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_742  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_743  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_744  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_745  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_746  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_747  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_748  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_749  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_750  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_751  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_752  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_753  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_754  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_755  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_756  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_757  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_758  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_759  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_760  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_761  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_762  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_763  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_764  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_765  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_766  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_767  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_768  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_769  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_770  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_771  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_772  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_773  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_774  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_775  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_776  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_777  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_778  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_779  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_780  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_781  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_782  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_783  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_784  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_785  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_786  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_787  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_788  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_789  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_790  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_791  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_792  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_793  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_794  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_795  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_796  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_797  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_798  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_799  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_800  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_801  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_802  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_803  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_804  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_805  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_806  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_807  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_808  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_809  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_810  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_811  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_812  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_813  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_814  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_815  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_816  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_817  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_818  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_819  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_820  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_821  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_822  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_823  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_824  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_825  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_826  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_827  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_828  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_829  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_830  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_831  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_832  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_833  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_834  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_835  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_836  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_837  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_838  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_839  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_840  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_841  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_842  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_843  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_844  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_845  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_846  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_847  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_848  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_849  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_850  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_851  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_852  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_853  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_854  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_855  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_856  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_857  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_858  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_859  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_860  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_861  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_862  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_863  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_864  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_865  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_866  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_867  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_868  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_869  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_870  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_871  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_872  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_873  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_874  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_875  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_876  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_877  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_878  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_879  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_880  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_881  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_882  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_883  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_884  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_885  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_886  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_887  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_888  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_889  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_890  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_891  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_892  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_893  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_894  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_895  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_896  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_897  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_898  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_899  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_900  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_901  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_902  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_903  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_904  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_905  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_906  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_907  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_908  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_909  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_910  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_911  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_912  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_913  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_914  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_915  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_916  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_917  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_918  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_919  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_920  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_921  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_922  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_923  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_924  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_925  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_926  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_927  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_928  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_929  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_930  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_931  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_932  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_933  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_934  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_935  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_936  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_937  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_938  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_939  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_940  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_941  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_942  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_943  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_944  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_945  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_946  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_947  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_948  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_949  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_950  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_951  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_952  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_953  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_954  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_955  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_956  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_957  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_958  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_959  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_960  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_961  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_962  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_963  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_964  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_965  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_966  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_967  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_968  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_969  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_970  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_971  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_972  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_973  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_974  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_975  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_976  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_977  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_978  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_979  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_980  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_981  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_982  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_983  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_984  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_985  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_986  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_987  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_988  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_989  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_990  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_991  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_992  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_993  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_994  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_995  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_996  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_997  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_998  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_999  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1000 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1001 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1002 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1003 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1004 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1005 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1006 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1007 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1008 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1009 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1010 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1011 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1012 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1013 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1014 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1015 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1016 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1017 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1018 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1019 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1020 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1021 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1022 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1023 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1024 :out std_logic_vector(11 downto 0)

       );

end component PeakDetector;

component TB_ReadAdc is
  --+----------
  -- Generic declarations
  --+----------
  generic(
          DataVecSize_g   :integer := 56;
          WdVecSize_g     :integer := 16;
          ByteSize_g      :integer := 8;
          NibbleSize_g    :integer := 4
      );

  --+----------
  -- Port name declarations
  --+----------
  port   (
       CLK100              :in  std_logic;
       RST                 :in  std_logic;
--       TEST              :in  std_logic;       
       ADC_CLK_1           :out std_logic;   
       ADC_CLK_2           :out std_logic;

       i_DR1_EN            :in std_logic;
       i_DR2_EN            :in std_logic;
       
       ADC_D1              :in  std_logic_vector(WdVecSize_g-5 downto 0);
       ADC_DR1             :in  std_logic;
       
       ADC_D2              :in  std_logic_vector(WdVecSize_g-5 downto 0);
       ADC_DR2             :in  std_logic;

       DATA1       :out std_logic_vector(WdVecSize_g-5 downto 0);
       DATARDY1    :out std_logic;
       
       DATA2       :out std_logic_vector(WdVecSize_g-5 downto 0);
       DATARDY2    :out std_logic;
	   
	   i_stop_req  :in  std_logic

         );

end component TB_ReadAdc;

--+----------
-- Start of architecture code
--+----------
begin
  --+----------
  -- Global signal assignments for the architecture.
  --+----------
-- STOP    <= Stop_s;

  i_reset_n  <= not RST;
 
 PEAK_FL_C1    <=  PEAK_FL_C1_s;

 PEAK_C1       <=  PEAK_C1_s;
--PEAK_C2       <=  PEAK_C2_s;

 ADC_D1_s      <=   ADC_D1_d;   
 ADC_DR1_s     <=   ADC_DR1_d;
 ADC_D2_s      <=   ADC_D2_d ;
 ADC_DR2_s     <=   ADC_DR2_d;
 
 --data_update_process : process(CLK100, RST)
 --begin
    --if(RST = '1') then
         --energy_bin_pos_data(954 ) <= (others=>'0');
    --elsif rising_edge(CLK100) then
        --energy_bin_pos_data(954 ) <= s_energy_bin_pos_data_954;
    --end if;
    --
 --end process data_update_process;
 
-- ************************************************************************************************************************ adc data fifos ******************************************************************************************************
adc_data_fifo_inst_1 : adc_data_fifo
port map(
        CLK     => CLK100,
        DATA    => adc_fifo_data_in_1,
        RE      => rd_en_adc_fifo_1,
        RESET_N => i_reset_n,
        WE      => wr_en_adc_fifo_1,
        EMPTY   => adc_fifo_empty_1,
        FULL    => adc_fifo_full_1,
        Q       => adc_fifo_data_out_1
);

adc_data_fifo_inst_2 : adc_data_fifo
port map(
        CLK     => CLK100,
        DATA    => adc_fifo_data_in_2,
        RE      => rd_en_adc_fifo_2,
        RESET_N => i_reset_n,
        WE      => wr_en_adc_fifo_2,
        EMPTY   => adc_fifo_empty_2,
        FULL    => adc_fifo_full_2,
        Q       => adc_fifo_data_out_2
);

--****************************************************************************************************peak data fifos****************************************************************************************************************************

peak_fifo_inst_1 : peak_data_fifo
port map(
        CLK     => CLK100,
        DATA    => peak_fifo_data_in_1,
        RE      => rd_en_peak_fifo_1,
        RESET_N => i_reset_n,
        WE      => wr_en_peak_fifo_1,
        EMPTY   => peak_fifo_empty_1,
        FULL    => peak_fifo_full_1,
        Q       => peak_fifo_data_out_1
);

peak_fifo_inst_2 : peak_data_fifo
port map(
        CLK     => CLK100,
        DATA    => peak_fifo_data_in_2,
        RE      => rd_en_peak_fifo_2,
        RESET_N => i_reset_n,
        WE      => wr_en_peak_fifo_2,
        EMPTY   => peak_fifo_empty_2,
        FULL    => peak_fifo_full_2,
        Q       => peak_fifo_data_out_2
);

TimeStampCtrl_inst : TimeStampCtrl

  port map  (
       CLK100        =>   CLK100,
       RST           =>   RST,
       DATARDY1      =>   DATARDY1,
       DATARDY2      =>   DATARDY2,
       TIMESTAMP_C1  =>   TIMESTAMP_C1,
       TIMESTAMP_C2  =>   TIMESTAMP_C2
         );

PeakDetector_inst :PeakDetector
  port map  (
       CLK100                =>   CLK100,
       RST                   =>   RST,
       
       DATA1                 =>   DATA1    ,
       DATARDY1              =>   DATARDY1 ,  
       DATA2                 =>   DATA2    ,
       DATARDY2              =>   DATARDY2 ,
       
       ADD_TIMP_FLAG  	     =>   PEAK_FL_C1_s ,    
       ADD_TIMP_FLAG_pos     =>   PEAK_FL_C1_s_pos ,    
       o_DATA_OUT_C1         =>   PEAK_C1_s    ,     
       o_DATA_OUT_C2         =>   PEAK_C1_s_pos    ,

	   o_Energy_Bin_Pos_1    =>   energy_bin_pos_data(0	  ),
	   o_Energy_Bin_Pos_2    =>   energy_bin_pos_data(1   ),
	   o_Energy_Bin_Pos_3    =>   energy_bin_pos_data(2   ),
	   o_Energy_Bin_Pos_4    =>   energy_bin_pos_data(3   ),
	   o_Energy_Bin_Pos_5    =>   energy_bin_pos_data(4   ),
	   o_Energy_Bin_Pos_6    =>   energy_bin_pos_data(5   ),
	   o_Energy_Bin_Pos_7    =>   energy_bin_pos_data(6   ),
	   o_Energy_Bin_Pos_8    =>   energy_bin_pos_data(7   ),
	   o_Energy_Bin_Pos_9    =>   energy_bin_pos_data(8   ),
	   o_Energy_Bin_Pos_10   =>   energy_bin_pos_data(9   ),
	   o_Energy_Bin_Pos_11   =>   energy_bin_pos_data(10  ),
	   o_Energy_Bin_Pos_12   =>   energy_bin_pos_data(11  ),
	   o_Energy_Bin_Pos_13   =>   energy_bin_pos_data(12  ),
	   o_Energy_Bin_Pos_14   =>   energy_bin_pos_data(13  ),
	   o_Energy_Bin_Pos_15   =>   energy_bin_pos_data(14  ),
	   o_Energy_Bin_Pos_16   =>   energy_bin_pos_data(15  ),
	   o_Energy_Bin_Pos_17   =>   energy_bin_pos_data(16  ),
	   o_Energy_Bin_Pos_18   =>   energy_bin_pos_data(17  ),
	   o_Energy_Bin_Pos_19   =>   energy_bin_pos_data(18  ),
	   o_Energy_Bin_Pos_20   =>   energy_bin_pos_data(19  ),
	   o_Energy_Bin_Pos_21   =>   energy_bin_pos_data(20  ),
	   o_Energy_Bin_Pos_22   =>   energy_bin_pos_data(21  ),
	   o_Energy_Bin_Pos_23   =>   energy_bin_pos_data(22  ),
	   o_Energy_Bin_Pos_24   =>   energy_bin_pos_data(23  ),
	   o_Energy_Bin_Pos_25   =>   energy_bin_pos_data(24  ),
	   o_Energy_Bin_Pos_26   =>   energy_bin_pos_data(25  ),
	   o_Energy_Bin_Pos_27   =>   energy_bin_pos_data(26  ),
	   o_Energy_Bin_Pos_28   =>   energy_bin_pos_data(27  ),
	   o_Energy_Bin_Pos_29   =>   energy_bin_pos_data(28  ),
	   o_Energy_Bin_Pos_30   =>   energy_bin_pos_data(29  ),
	   o_Energy_Bin_Pos_31   =>   energy_bin_pos_data(30  ),
	   o_Energy_Bin_Pos_32   =>   energy_bin_pos_data(31  ),
	   o_Energy_Bin_Pos_33   =>   energy_bin_pos_data(32  ),
	   o_Energy_Bin_Pos_34   =>   energy_bin_pos_data(33  ),
	   o_Energy_Bin_Pos_35   =>   energy_bin_pos_data(34  ),
	   o_Energy_Bin_Pos_36   =>   energy_bin_pos_data(35  ),
	   o_Energy_Bin_Pos_37   =>   energy_bin_pos_data(36  ),
	   o_Energy_Bin_Pos_38   =>   energy_bin_pos_data(37  ),
	   o_Energy_Bin_Pos_39   =>   energy_bin_pos_data(38  ),
	   o_Energy_Bin_Pos_40   =>   energy_bin_pos_data(39  ),
	   o_Energy_Bin_Pos_41   =>   energy_bin_pos_data(40  ),
	   o_Energy_Bin_Pos_42   =>   energy_bin_pos_data(41  ),
	   o_Energy_Bin_Pos_43   =>   energy_bin_pos_data(42  ),
	   o_Energy_Bin_Pos_44   =>   energy_bin_pos_data(43  ),
	   o_Energy_Bin_Pos_45   =>   energy_bin_pos_data(44  ),
	   o_Energy_Bin_Pos_46   =>   energy_bin_pos_data(45  ),
	   o_Energy_Bin_Pos_47   =>   energy_bin_pos_data(46  ),
	   o_Energy_Bin_Pos_48   =>   energy_bin_pos_data(47  ),
	   o_Energy_Bin_Pos_49   =>   energy_bin_pos_data(48  ),
	   o_Energy_Bin_Pos_50   =>   energy_bin_pos_data(49  ),
	   o_Energy_Bin_Pos_51   =>   energy_bin_pos_data(50  ),
	   o_Energy_Bin_Pos_52   =>   energy_bin_pos_data(51  ),
	   o_Energy_Bin_Pos_53   =>   energy_bin_pos_data(52  ),
	   o_Energy_Bin_Pos_54   =>   energy_bin_pos_data(53  ),
	   o_Energy_Bin_Pos_55   =>   energy_bin_pos_data(54  ),
	   o_Energy_Bin_Pos_56   =>   energy_bin_pos_data(55  ),
	   o_Energy_Bin_Pos_57   =>   energy_bin_pos_data(56  ),
	   o_Energy_Bin_Pos_58   =>   energy_bin_pos_data(57  ),
	   o_Energy_Bin_Pos_59   =>   energy_bin_pos_data(58  ),
	   o_Energy_Bin_Pos_60   =>   energy_bin_pos_data(59  ),
	   o_Energy_Bin_Pos_61   =>   energy_bin_pos_data(60  ),
	   o_Energy_Bin_Pos_62   =>   energy_bin_pos_data(61  ),
	   o_Energy_Bin_Pos_63   =>   energy_bin_pos_data(62  ),
	   o_Energy_Bin_Pos_64   =>   energy_bin_pos_data(63  ),
	   o_Energy_Bin_Pos_65   =>   energy_bin_pos_data(64  ),
	   o_Energy_Bin_Pos_66   =>   energy_bin_pos_data(65  ),
	   o_Energy_Bin_Pos_67   =>   energy_bin_pos_data(66  ),
	   o_Energy_Bin_Pos_68   =>   energy_bin_pos_data(67  ),
	   o_Energy_Bin_Pos_69   =>   energy_bin_pos_data(68  ),
	   o_Energy_Bin_Pos_70   =>   energy_bin_pos_data(69  ),
	   o_Energy_Bin_Pos_71   =>   energy_bin_pos_data(70  ),
	   o_Energy_Bin_Pos_72   =>   energy_bin_pos_data(71  ),
	   o_Energy_Bin_Pos_73   =>   energy_bin_pos_data(72  ),
	   o_Energy_Bin_Pos_74   =>   energy_bin_pos_data(73  ),
	   o_Energy_Bin_Pos_75   =>   energy_bin_pos_data(74  ),
	   o_Energy_Bin_Pos_76   =>   energy_bin_pos_data(75  ),
	   o_Energy_Bin_Pos_77   =>   energy_bin_pos_data(76  ),
	   o_Energy_Bin_Pos_78   =>   energy_bin_pos_data(77  ),
	   o_Energy_Bin_Pos_79   =>   energy_bin_pos_data(78  ),
	   o_Energy_Bin_Pos_80   =>   energy_bin_pos_data(79  ),
	   o_Energy_Bin_Pos_81   =>   energy_bin_pos_data(80  ),
	   o_Energy_Bin_Pos_82   =>   energy_bin_pos_data(81  ),
	   o_Energy_Bin_Pos_83   =>   energy_bin_pos_data(82  ),
	   o_Energy_Bin_Pos_84   =>   energy_bin_pos_data(83  ),
	   o_Energy_Bin_Pos_85   =>   energy_bin_pos_data(84  ),
	   o_Energy_Bin_Pos_86   =>   energy_bin_pos_data(85  ),
	   o_Energy_Bin_Pos_87   =>   energy_bin_pos_data(86  ),
	   o_Energy_Bin_Pos_88   =>   energy_bin_pos_data(87  ),
	   o_Energy_Bin_Pos_89   =>   energy_bin_pos_data(88  ),
	   o_Energy_Bin_Pos_90   =>   energy_bin_pos_data(89  ),
	   o_Energy_Bin_Pos_91   =>   energy_bin_pos_data(90  ),
	   o_Energy_Bin_Pos_92   =>   energy_bin_pos_data(91  ),
	   o_Energy_Bin_Pos_93   =>   energy_bin_pos_data(92  ),
	   o_Energy_Bin_Pos_94   =>   energy_bin_pos_data(93  ),
	   o_Energy_Bin_Pos_95   =>   energy_bin_pos_data(94  ),
	   o_Energy_Bin_Pos_96   =>   energy_bin_pos_data(95  ),
	   o_Energy_Bin_Pos_97   =>   energy_bin_pos_data(96  ),
	   o_Energy_Bin_Pos_98   =>   energy_bin_pos_data(97  ),
	   o_Energy_Bin_Pos_99   =>   energy_bin_pos_data(98  ),
	   o_Energy_Bin_Pos_100  =>   energy_bin_pos_data(99  ),
	   o_Energy_Bin_Pos_101  =>   energy_bin_pos_data(100 ),
	   o_Energy_Bin_Pos_102  =>   energy_bin_pos_data(101 ),
	   o_Energy_Bin_Pos_103  =>   energy_bin_pos_data(102 ),
	   o_Energy_Bin_Pos_104  =>   energy_bin_pos_data(103 ),
	   o_Energy_Bin_Pos_105  =>   energy_bin_pos_data(104 ),
	   o_Energy_Bin_Pos_106  =>   energy_bin_pos_data(105 ),
	   o_Energy_Bin_Pos_107  =>   energy_bin_pos_data(106 ),
	   o_Energy_Bin_Pos_108  =>   energy_bin_pos_data(107 ),
	   o_Energy_Bin_Pos_109  =>   energy_bin_pos_data(108 ),
	   o_Energy_Bin_Pos_110  =>   energy_bin_pos_data(109 ),
	   o_Energy_Bin_Pos_111  =>   energy_bin_pos_data(110 ),
	   o_Energy_Bin_Pos_112  =>   energy_bin_pos_data(111 ),
	   o_Energy_Bin_Pos_113  =>   energy_bin_pos_data(112 ),
	   o_Energy_Bin_Pos_114  =>   energy_bin_pos_data(113 ),
	   o_Energy_Bin_Pos_115  =>   energy_bin_pos_data(114 ),
	   o_Energy_Bin_Pos_116  =>   energy_bin_pos_data(115 ),
	   o_Energy_Bin_Pos_117  =>   energy_bin_pos_data(116 ),
	   o_Energy_Bin_Pos_118  =>   energy_bin_pos_data(117 ),
	   o_Energy_Bin_Pos_119  =>   energy_bin_pos_data(118 ),
	   o_Energy_Bin_Pos_120  =>   energy_bin_pos_data(119 ),
	   o_Energy_Bin_Pos_121  =>   energy_bin_pos_data(120 ),
	   o_Energy_Bin_Pos_122  =>   energy_bin_pos_data(121 ),
	   o_Energy_Bin_Pos_123  =>   energy_bin_pos_data(122 ),
	   o_Energy_Bin_Pos_124  =>   energy_bin_pos_data(123 ),
	   o_Energy_Bin_Pos_125  =>   energy_bin_pos_data(124 ),
	   o_Energy_Bin_Pos_126  =>   energy_bin_pos_data(125 ),
	   o_Energy_Bin_Pos_127  =>   energy_bin_pos_data(126 ),
	   o_Energy_Bin_Pos_128  =>   energy_bin_pos_data(127 ),
	   o_Energy_Bin_Pos_129  =>   energy_bin_pos_data(128 ),
	   o_Energy_Bin_Pos_130  =>   energy_bin_pos_data(129 ),
	   o_Energy_Bin_Pos_131  =>   energy_bin_pos_data(130 ),
	   o_Energy_Bin_Pos_132  =>   energy_bin_pos_data(131 ),
	   o_Energy_Bin_Pos_133  =>   energy_bin_pos_data(132 ),
	   o_Energy_Bin_Pos_134  =>   energy_bin_pos_data(133 ),
	   o_Energy_Bin_Pos_135  =>   energy_bin_pos_data(134 ),
	   o_Energy_Bin_Pos_136  =>   energy_bin_pos_data(135 ),
	   o_Energy_Bin_Pos_137  =>   energy_bin_pos_data(136 ),
	   o_Energy_Bin_Pos_138  =>   energy_bin_pos_data(137 ),
	   o_Energy_Bin_Pos_139  =>   energy_bin_pos_data(138 ),
	   o_Energy_Bin_Pos_140  =>   energy_bin_pos_data(139 ),
	   o_Energy_Bin_Pos_141  =>   energy_bin_pos_data(140 ),
	   o_Energy_Bin_Pos_142  =>   energy_bin_pos_data(141 ),
	   o_Energy_Bin_Pos_143  =>   energy_bin_pos_data(142 ),
	   o_Energy_Bin_Pos_144  =>   energy_bin_pos_data(143 ),
	   o_Energy_Bin_Pos_145  =>   energy_bin_pos_data(144 ),
	   o_Energy_Bin_Pos_146  =>   energy_bin_pos_data(145 ),
	   o_Energy_Bin_Pos_147  =>   energy_bin_pos_data(146 ),
	   o_Energy_Bin_Pos_148  =>   energy_bin_pos_data(147 ),
	   o_Energy_Bin_Pos_149  =>   energy_bin_pos_data(148 ),
	   o_Energy_Bin_Pos_150  =>   energy_bin_pos_data(149 ),
	   o_Energy_Bin_Pos_151  =>   energy_bin_pos_data(150 ),
	   o_Energy_Bin_Pos_152  =>   energy_bin_pos_data(151 ),
	   o_Energy_Bin_Pos_153  =>   energy_bin_pos_data(152 ),
	   o_Energy_Bin_Pos_154  =>   energy_bin_pos_data(153 ),
	   o_Energy_Bin_Pos_155  =>   energy_bin_pos_data(154 ),
	   o_Energy_Bin_Pos_156  =>   energy_bin_pos_data(155 ),
	   o_Energy_Bin_Pos_157  =>   energy_bin_pos_data(156 ),
	   o_Energy_Bin_Pos_158  =>   energy_bin_pos_data(157 ),
	   o_Energy_Bin_Pos_159  =>   energy_bin_pos_data(158 ),
	   o_Energy_Bin_Pos_160  =>   energy_bin_pos_data(159 ),
	   o_Energy_Bin_Pos_161  =>   energy_bin_pos_data(160 ),
	   o_Energy_Bin_Pos_162  =>   energy_bin_pos_data(161 ),
	   o_Energy_Bin_Pos_163  =>   energy_bin_pos_data(162 ),
	   o_Energy_Bin_Pos_164  =>   energy_bin_pos_data(163 ),
	   o_Energy_Bin_Pos_165  =>   energy_bin_pos_data(164 ),
	   o_Energy_Bin_Pos_166  =>   energy_bin_pos_data(165 ),
	   o_Energy_Bin_Pos_167  =>   energy_bin_pos_data(166 ),
	   o_Energy_Bin_Pos_168  =>   energy_bin_pos_data(167 ),
	   o_Energy_Bin_Pos_169  =>   energy_bin_pos_data(168 ),
	   o_Energy_Bin_Pos_170  =>   energy_bin_pos_data(169 ),
	   o_Energy_Bin_Pos_171  =>   energy_bin_pos_data(170 ),
	   o_Energy_Bin_Pos_172  =>   energy_bin_pos_data(171 ),
	   o_Energy_Bin_Pos_173  =>   energy_bin_pos_data(172 ),
	   o_Energy_Bin_Pos_174  =>   energy_bin_pos_data(173 ),
	   o_Energy_Bin_Pos_175  =>   energy_bin_pos_data(174 ),
	   o_Energy_Bin_Pos_176  =>   energy_bin_pos_data(175 ),
	   o_Energy_Bin_Pos_177  =>   energy_bin_pos_data(176 ),
	   o_Energy_Bin_Pos_178  =>   energy_bin_pos_data(177 ),
	   o_Energy_Bin_Pos_179  =>   energy_bin_pos_data(178 ),
	   o_Energy_Bin_Pos_180  =>   energy_bin_pos_data(179 ),
	   o_Energy_Bin_Pos_181  =>   energy_bin_pos_data(180 ),
	   o_Energy_Bin_Pos_182  =>   energy_bin_pos_data(181 ),
	   o_Energy_Bin_Pos_183  =>   energy_bin_pos_data(182 ),
	   o_Energy_Bin_Pos_184  =>   energy_bin_pos_data(183 ),
	   o_Energy_Bin_Pos_185  =>   energy_bin_pos_data(184 ),
	   o_Energy_Bin_Pos_186  =>   energy_bin_pos_data(185 ),
	   o_Energy_Bin_Pos_187  =>   energy_bin_pos_data(186 ),
	   o_Energy_Bin_Pos_188  =>   energy_bin_pos_data(187 ),
	   o_Energy_Bin_Pos_189  =>   energy_bin_pos_data(188 ),
	   o_Energy_Bin_Pos_190  =>   energy_bin_pos_data(189 ),
	   o_Energy_Bin_Pos_191  =>   energy_bin_pos_data(190 ),
	   o_Energy_Bin_Pos_192  =>   energy_bin_pos_data(191 ),
	   o_Energy_Bin_Pos_193  =>   energy_bin_pos_data(192 ),
	   o_Energy_Bin_Pos_194  =>   energy_bin_pos_data(193 ),
	   o_Energy_Bin_Pos_195  =>   energy_bin_pos_data(194 ),
	   o_Energy_Bin_Pos_196  =>   energy_bin_pos_data(195 ),
	   o_Energy_Bin_Pos_197  =>   energy_bin_pos_data(196 ),
	   o_Energy_Bin_Pos_198  =>   energy_bin_pos_data(197 ),
	   o_Energy_Bin_Pos_199  =>   energy_bin_pos_data(198 ),
	   o_Energy_Bin_Pos_200  =>   energy_bin_pos_data(199 ),
	   o_Energy_Bin_Pos_201  =>   energy_bin_pos_data(200 ),
	   o_Energy_Bin_Pos_202  =>   energy_bin_pos_data(201 ),
	   o_Energy_Bin_Pos_203  =>   energy_bin_pos_data(202 ),
	   o_Energy_Bin_Pos_204  =>   energy_bin_pos_data(203 ),
	   o_Energy_Bin_Pos_205  =>   energy_bin_pos_data(204 ),
	   o_Energy_Bin_Pos_206  =>   energy_bin_pos_data(205 ),
	   o_Energy_Bin_Pos_207  =>   energy_bin_pos_data(206 ),
	   o_Energy_Bin_Pos_208  =>   energy_bin_pos_data(207 ),
	   o_Energy_Bin_Pos_209  =>   energy_bin_pos_data(208 ),
	   o_Energy_Bin_Pos_210  =>   energy_bin_pos_data(209 ),
	   o_Energy_Bin_Pos_211  =>   energy_bin_pos_data(210 ),
	   o_Energy_Bin_Pos_212  =>   energy_bin_pos_data(211 ),
	   o_Energy_Bin_Pos_213  =>   energy_bin_pos_data(212 ),
	   o_Energy_Bin_Pos_214  =>   energy_bin_pos_data(213 ),
	   o_Energy_Bin_Pos_215  =>   energy_bin_pos_data(214 ),
	   o_Energy_Bin_Pos_216  =>   energy_bin_pos_data(215 ),
	   o_Energy_Bin_Pos_217  =>   energy_bin_pos_data(216 ),
	   o_Energy_Bin_Pos_218  =>   energy_bin_pos_data(217 ),
	   o_Energy_Bin_Pos_219  =>   energy_bin_pos_data(218 ),
	   o_Energy_Bin_Pos_220  =>   energy_bin_pos_data(219 ),
	   o_Energy_Bin_Pos_221  =>   energy_bin_pos_data(220 ),
	   o_Energy_Bin_Pos_222  =>   energy_bin_pos_data(221 ),
	   o_Energy_Bin_Pos_223  =>   energy_bin_pos_data(222 ),
	   o_Energy_Bin_Pos_224  =>   energy_bin_pos_data(223 ),
	   o_Energy_Bin_Pos_225  =>   energy_bin_pos_data(224 ),
	   o_Energy_Bin_Pos_226  =>   energy_bin_pos_data(225 ),
	   o_Energy_Bin_Pos_227  =>   energy_bin_pos_data(226 ),
	   o_Energy_Bin_Pos_228  =>   energy_bin_pos_data(227 ),
	   o_Energy_Bin_Pos_229  =>   energy_bin_pos_data(228 ),
	   o_Energy_Bin_Pos_230  =>   energy_bin_pos_data(229 ),
	   o_Energy_Bin_Pos_231  =>   energy_bin_pos_data(230 ),
	   o_Energy_Bin_Pos_232  =>   energy_bin_pos_data(231 ),
	   o_Energy_Bin_Pos_233  =>   energy_bin_pos_data(232 ),
	   o_Energy_Bin_Pos_234  =>   energy_bin_pos_data(233 ),
	   o_Energy_Bin_Pos_235  =>   energy_bin_pos_data(234 ),
	   o_Energy_Bin_Pos_236  =>   energy_bin_pos_data(235 ),
	   o_Energy_Bin_Pos_237  =>   energy_bin_pos_data(236 ),
	   o_Energy_Bin_Pos_238  =>   energy_bin_pos_data(237 ),
	   o_Energy_Bin_Pos_239  =>   energy_bin_pos_data(238 ),
	   o_Energy_Bin_Pos_240  =>   energy_bin_pos_data(239 ),
	   o_Energy_Bin_Pos_241  =>   energy_bin_pos_data(240 ),
	   o_Energy_Bin_Pos_242  =>   energy_bin_pos_data(241 ),
	   o_Energy_Bin_Pos_243  =>   energy_bin_pos_data(242 ),
	   o_Energy_Bin_Pos_244  =>   energy_bin_pos_data(243 ),
	   o_Energy_Bin_Pos_245  =>   energy_bin_pos_data(244 ),
	   o_Energy_Bin_Pos_246  =>   energy_bin_pos_data(245 ),
	   o_Energy_Bin_Pos_247  =>   energy_bin_pos_data(246 ),
	   o_Energy_Bin_Pos_248  =>   energy_bin_pos_data(247 ),
	   o_Energy_Bin_Pos_249  =>   energy_bin_pos_data(248 ),
	   o_Energy_Bin_Pos_250  =>   energy_bin_pos_data(249 ),
	   o_Energy_Bin_Pos_251  =>   energy_bin_pos_data(250 ),
	   o_Energy_Bin_Pos_252  =>   energy_bin_pos_data(251 ),
	   o_Energy_Bin_Pos_253  =>   energy_bin_pos_data(252 ),
	   o_Energy_Bin_Pos_254  =>   energy_bin_pos_data(253 ),
	   o_Energy_Bin_Pos_255  =>   energy_bin_pos_data(254 ),
	   o_Energy_Bin_Pos_256  =>   energy_bin_pos_data(255 ),
	   o_Energy_Bin_Pos_257  =>   energy_bin_pos_data(256 ),
	   o_Energy_Bin_Pos_258  =>   energy_bin_pos_data(257 ),
	   o_Energy_Bin_Pos_259  =>   energy_bin_pos_data(258 ),
	   o_Energy_Bin_Pos_260  =>   energy_bin_pos_data(259 ),
	   o_Energy_Bin_Pos_261  =>   energy_bin_pos_data(260 ),
	   o_Energy_Bin_Pos_262  =>   energy_bin_pos_data(261 ),
	   o_Energy_Bin_Pos_263  =>   energy_bin_pos_data(262 ),
	   o_Energy_Bin_Pos_264  =>   energy_bin_pos_data(263 ),
	   o_Energy_Bin_Pos_265  =>   energy_bin_pos_data(264 ),
	   o_Energy_Bin_Pos_266  =>   energy_bin_pos_data(265 ),
	   o_Energy_Bin_Pos_267  =>   energy_bin_pos_data(266 ),
	   o_Energy_Bin_Pos_268  =>   energy_bin_pos_data(267 ),
	   o_Energy_Bin_Pos_269  =>   energy_bin_pos_data(268 ),
	   o_Energy_Bin_Pos_270  =>   energy_bin_pos_data(269 ),
	   o_Energy_Bin_Pos_271  =>   energy_bin_pos_data(270 ),
	   o_Energy_Bin_Pos_272  =>   energy_bin_pos_data(271 ),
	   o_Energy_Bin_Pos_273  =>   energy_bin_pos_data(272 ),
	   o_Energy_Bin_Pos_274  =>   energy_bin_pos_data(273 ),
	   o_Energy_Bin_Pos_275  =>   energy_bin_pos_data(274 ),
	   o_Energy_Bin_Pos_276  =>   energy_bin_pos_data(275 ),
	   o_Energy_Bin_Pos_277  =>   energy_bin_pos_data(276 ),
	   o_Energy_Bin_Pos_278  =>   energy_bin_pos_data(277 ),
	   o_Energy_Bin_Pos_279  =>   energy_bin_pos_data(278 ),
	   o_Energy_Bin_Pos_280  =>   energy_bin_pos_data(279 ),
	   o_Energy_Bin_Pos_281  =>   energy_bin_pos_data(280 ),
	   o_Energy_Bin_Pos_282  =>   energy_bin_pos_data(281 ),
	   o_Energy_Bin_Pos_283  =>   energy_bin_pos_data(282 ),
	   o_Energy_Bin_Pos_284  =>   energy_bin_pos_data(283 ),
	   o_Energy_Bin_Pos_285  =>   energy_bin_pos_data(284 ),
	   o_Energy_Bin_Pos_286  =>   energy_bin_pos_data(285 ),
	   o_Energy_Bin_Pos_287  =>   energy_bin_pos_data(286 ),
	   o_Energy_Bin_Pos_288  =>   energy_bin_pos_data(287 ),
	   o_Energy_Bin_Pos_289  =>   energy_bin_pos_data(288 ),
	   o_Energy_Bin_Pos_290  =>   energy_bin_pos_data(289 ),
	   o_Energy_Bin_Pos_291  =>   energy_bin_pos_data(290 ),
	   o_Energy_Bin_Pos_292  =>   energy_bin_pos_data(291 ),
	   o_Energy_Bin_Pos_293  =>   energy_bin_pos_data(292 ),
	   o_Energy_Bin_Pos_294  =>   energy_bin_pos_data(293 ),
	   o_Energy_Bin_Pos_295  =>   energy_bin_pos_data(294 ),
	   o_Energy_Bin_Pos_296  =>   energy_bin_pos_data(295 ),
	   o_Energy_Bin_Pos_297  =>   energy_bin_pos_data(296 ),
	   o_Energy_Bin_Pos_298  =>   energy_bin_pos_data(297 ),
	   o_Energy_Bin_Pos_299  =>   energy_bin_pos_data(298 ),
	   o_Energy_Bin_Pos_300  =>   energy_bin_pos_data(299 ),
	   o_Energy_Bin_Pos_301  =>   energy_bin_pos_data(300 ),
	   o_Energy_Bin_Pos_302  =>   energy_bin_pos_data(301 ),
	   o_Energy_Bin_Pos_303  =>   energy_bin_pos_data(302 ),
	   o_Energy_Bin_Pos_304  =>   energy_bin_pos_data(303 ),
	   o_Energy_Bin_Pos_305  =>   energy_bin_pos_data(304 ),
	   o_Energy_Bin_Pos_306  =>   energy_bin_pos_data(305 ),
	   o_Energy_Bin_Pos_307  =>   energy_bin_pos_data(306 ),
	   o_Energy_Bin_Pos_308  =>   energy_bin_pos_data(307 ),
	   o_Energy_Bin_Pos_309  =>   energy_bin_pos_data(308 ),
	   o_Energy_Bin_Pos_310  =>   energy_bin_pos_data(309 ),
	   o_Energy_Bin_Pos_311  =>   energy_bin_pos_data(310 ),
	   o_Energy_Bin_Pos_312  =>   energy_bin_pos_data(311 ),
	   o_Energy_Bin_Pos_313  =>   energy_bin_pos_data(312 ),
	   o_Energy_Bin_Pos_314  =>   energy_bin_pos_data(313 ),
	   o_Energy_Bin_Pos_315  =>   energy_bin_pos_data(314 ),
	   o_Energy_Bin_Pos_316  =>   energy_bin_pos_data(315 ),
	   o_Energy_Bin_Pos_317  =>   energy_bin_pos_data(316 ),
	   o_Energy_Bin_Pos_318  =>   energy_bin_pos_data(317 ),
	   o_Energy_Bin_Pos_319  =>   energy_bin_pos_data(318 ),
	   o_Energy_Bin_Pos_320  =>   energy_bin_pos_data(319 ),
	   o_Energy_Bin_Pos_321  =>   energy_bin_pos_data(320 ),
	   o_Energy_Bin_Pos_322  =>   energy_bin_pos_data(321 ),
	   o_Energy_Bin_Pos_323  =>   energy_bin_pos_data(322 ),
	   o_Energy_Bin_Pos_324  =>   energy_bin_pos_data(323 ),
	   o_Energy_Bin_Pos_325  =>   energy_bin_pos_data(324 ),
	   o_Energy_Bin_Pos_326  =>   energy_bin_pos_data(325 ),
	   o_Energy_Bin_Pos_327  =>   energy_bin_pos_data(326 ),
	   o_Energy_Bin_Pos_328  =>   energy_bin_pos_data(327 ),
	   o_Energy_Bin_Pos_329  =>   energy_bin_pos_data(328 ),
	   o_Energy_Bin_Pos_330  =>   energy_bin_pos_data(329 ),
	   o_Energy_Bin_Pos_331  =>   energy_bin_pos_data(330 ),
	   o_Energy_Bin_Pos_332  =>   energy_bin_pos_data(331 ),
	   o_Energy_Bin_Pos_333  =>   energy_bin_pos_data(332 ),
	   o_Energy_Bin_Pos_334  =>   energy_bin_pos_data(333 ),
	   o_Energy_Bin_Pos_335  =>   energy_bin_pos_data(334 ),
	   o_Energy_Bin_Pos_336  =>   energy_bin_pos_data(335 ),
	   o_Energy_Bin_Pos_337  =>   energy_bin_pos_data(336 ),
	   o_Energy_Bin_Pos_338  =>   energy_bin_pos_data(337 ),
	   o_Energy_Bin_Pos_339  =>   energy_bin_pos_data(338 ),
	   o_Energy_Bin_Pos_340  =>   energy_bin_pos_data(339 ),
	   o_Energy_Bin_Pos_341  =>   energy_bin_pos_data(340 ),
	   o_Energy_Bin_Pos_342  =>   energy_bin_pos_data(341 ),
	   o_Energy_Bin_Pos_343  =>   energy_bin_pos_data(342 ),
	   o_Energy_Bin_Pos_344  =>   energy_bin_pos_data(343 ),
	   o_Energy_Bin_Pos_345  =>   energy_bin_pos_data(344 ),
	   o_Energy_Bin_Pos_346  =>   energy_bin_pos_data(345 ),
	   o_Energy_Bin_Pos_347  =>   energy_bin_pos_data(346 ),
	   o_Energy_Bin_Pos_348  =>   energy_bin_pos_data(347 ),
	   o_Energy_Bin_Pos_349  =>   energy_bin_pos_data(348 ),
	   o_Energy_Bin_Pos_350  =>   energy_bin_pos_data(349 ),
	   o_Energy_Bin_Pos_351  =>   energy_bin_pos_data(350 ),
	   o_Energy_Bin_Pos_352  =>   energy_bin_pos_data(351 ),
	   o_Energy_Bin_Pos_353  =>   energy_bin_pos_data(352 ),
	   o_Energy_Bin_Pos_354  =>   energy_bin_pos_data(353 ),
	   o_Energy_Bin_Pos_355  =>   energy_bin_pos_data(354 ),
	   o_Energy_Bin_Pos_356  =>   energy_bin_pos_data(355 ),
	   o_Energy_Bin_Pos_357  =>   energy_bin_pos_data(356 ),
	   o_Energy_Bin_Pos_358  =>   energy_bin_pos_data(357 ),
	   o_Energy_Bin_Pos_359  =>   energy_bin_pos_data(358 ),
	   o_Energy_Bin_Pos_360  =>   energy_bin_pos_data(359 ),
	   o_Energy_Bin_Pos_361  =>   energy_bin_pos_data(360 ),
	   o_Energy_Bin_Pos_362  =>   energy_bin_pos_data(361 ),
	   o_Energy_Bin_Pos_363  =>   energy_bin_pos_data(362 ),
	   o_Energy_Bin_Pos_364  =>   energy_bin_pos_data(363 ),
	   o_Energy_Bin_Pos_365  =>   energy_bin_pos_data(364 ),
	   o_Energy_Bin_Pos_366  =>   energy_bin_pos_data(365 ),
	   o_Energy_Bin_Pos_367  =>   energy_bin_pos_data(366 ),
	   o_Energy_Bin_Pos_368  =>   energy_bin_pos_data(367 ),
	   o_Energy_Bin_Pos_369  =>   energy_bin_pos_data(368 ),
	   o_Energy_Bin_Pos_370  =>   energy_bin_pos_data(369 ),
	   o_Energy_Bin_Pos_371  =>   energy_bin_pos_data(370 ),
	   o_Energy_Bin_Pos_372  =>   energy_bin_pos_data(371 ),
	   o_Energy_Bin_Pos_373  =>   energy_bin_pos_data(372 ),
	   o_Energy_Bin_Pos_374  =>   energy_bin_pos_data(373 ),
	   o_Energy_Bin_Pos_375  =>   energy_bin_pos_data(374 ),
	   o_Energy_Bin_Pos_376  =>   energy_bin_pos_data(375 ),
	   o_Energy_Bin_Pos_377  =>   energy_bin_pos_data(376 ),
	   o_Energy_Bin_Pos_378  =>   energy_bin_pos_data(377 ),
	   o_Energy_Bin_Pos_379  =>   energy_bin_pos_data(378 ),
	   o_Energy_Bin_Pos_380  =>   energy_bin_pos_data(379 ),
	   o_Energy_Bin_Pos_381  =>   energy_bin_pos_data(380 ),
	   o_Energy_Bin_Pos_382  =>   energy_bin_pos_data(381 ),
	   o_Energy_Bin_Pos_383  =>   energy_bin_pos_data(382 ),
	   o_Energy_Bin_Pos_384  =>   energy_bin_pos_data(383 ),
	   o_Energy_Bin_Pos_385  =>   energy_bin_pos_data(384 ),
	   o_Energy_Bin_Pos_386  =>   energy_bin_pos_data(385 ),
	   o_Energy_Bin_Pos_387  =>   energy_bin_pos_data(386 ),
	   o_Energy_Bin_Pos_388  =>   energy_bin_pos_data(387 ),
	   o_Energy_Bin_Pos_389  =>   energy_bin_pos_data(388 ),
	   o_Energy_Bin_Pos_390  =>   energy_bin_pos_data(389 ),
	   o_Energy_Bin_Pos_391  =>   energy_bin_pos_data(390 ),
	   o_Energy_Bin_Pos_392  =>   energy_bin_pos_data(391 ),
	   o_Energy_Bin_Pos_393  =>   energy_bin_pos_data(392 ),
	   o_Energy_Bin_Pos_394  =>   energy_bin_pos_data(393 ),
	   o_Energy_Bin_Pos_395  =>   energy_bin_pos_data(394 ),
	   o_Energy_Bin_Pos_396  =>   energy_bin_pos_data(395 ),
	   o_Energy_Bin_Pos_397  =>   energy_bin_pos_data(396 ),
	   o_Energy_Bin_Pos_398  =>   energy_bin_pos_data(397 ),
	   o_Energy_Bin_Pos_399  =>   energy_bin_pos_data(398 ),
	   o_Energy_Bin_Pos_400  =>   energy_bin_pos_data(399 ),
	   o_Energy_Bin_Pos_401  =>   energy_bin_pos_data(400 ),
	   o_Energy_Bin_Pos_402  =>   energy_bin_pos_data(401 ),
	   o_Energy_Bin_Pos_403  =>   energy_bin_pos_data(402 ),
	   o_Energy_Bin_Pos_404  =>   energy_bin_pos_data(403 ),
	   o_Energy_Bin_Pos_405  =>   energy_bin_pos_data(404 ),
	   o_Energy_Bin_Pos_406  =>   energy_bin_pos_data(405 ),
	   o_Energy_Bin_Pos_407  =>   energy_bin_pos_data(406 ),
	   o_Energy_Bin_Pos_408  =>   energy_bin_pos_data(407 ),
	   o_Energy_Bin_Pos_409  =>   energy_bin_pos_data(408 ),
	   o_Energy_Bin_Pos_410  =>   energy_bin_pos_data(409 ),
	   o_Energy_Bin_Pos_411  =>   energy_bin_pos_data(410 ),
	   o_Energy_Bin_Pos_412  =>   energy_bin_pos_data(411 ),
	   o_Energy_Bin_Pos_413  =>   energy_bin_pos_data(412 ),
	   o_Energy_Bin_Pos_414  =>   energy_bin_pos_data(413 ),
	   o_Energy_Bin_Pos_415  =>   energy_bin_pos_data(414 ),
	   o_Energy_Bin_Pos_416  =>   energy_bin_pos_data(415 ),
	   o_Energy_Bin_Pos_417  =>   energy_bin_pos_data(416 ),
	   o_Energy_Bin_Pos_418  =>   energy_bin_pos_data(417 ),
	   o_Energy_Bin_Pos_419  =>   energy_bin_pos_data(418 ),
	   o_Energy_Bin_Pos_420  =>   energy_bin_pos_data(419 ),
	   o_Energy_Bin_Pos_421  =>   energy_bin_pos_data(420 ),
	   o_Energy_Bin_Pos_422  =>   energy_bin_pos_data(421 ),
	   o_Energy_Bin_Pos_423  =>   energy_bin_pos_data(422 ),
	   o_Energy_Bin_Pos_424  =>   energy_bin_pos_data(423 ),
	   o_Energy_Bin_Pos_425  =>   energy_bin_pos_data(424 ),
	   o_Energy_Bin_Pos_426  =>   energy_bin_pos_data(425 ),
	   o_Energy_Bin_Pos_427  =>   energy_bin_pos_data(426 ),
	   o_Energy_Bin_Pos_428  =>   energy_bin_pos_data(427 ),
	   o_Energy_Bin_Pos_429  =>   energy_bin_pos_data(428 ),
	   o_Energy_Bin_Pos_430  =>   energy_bin_pos_data(429 ),
	   o_Energy_Bin_Pos_431  =>   energy_bin_pos_data(430 ),
	   o_Energy_Bin_Pos_432  =>   energy_bin_pos_data(431 ),
	   o_Energy_Bin_Pos_433  =>   energy_bin_pos_data(432 ),
	   o_Energy_Bin_Pos_434  =>   energy_bin_pos_data(433 ),
	   o_Energy_Bin_Pos_435  =>   energy_bin_pos_data(434 ),
	   o_Energy_Bin_Pos_436  =>   energy_bin_pos_data(435 ),
	   o_Energy_Bin_Pos_437  =>   energy_bin_pos_data(436 ),
	   o_Energy_Bin_Pos_438  =>   energy_bin_pos_data(437 ),
	   o_Energy_Bin_Pos_439  =>   energy_bin_pos_data(438 ),
	   o_Energy_Bin_Pos_440  =>   energy_bin_pos_data(439 ),
	   o_Energy_Bin_Pos_441  =>   energy_bin_pos_data(440 ),
	   o_Energy_Bin_Pos_442  =>   energy_bin_pos_data(441 ),
	   o_Energy_Bin_Pos_443  =>   energy_bin_pos_data(442 ),
	   o_Energy_Bin_Pos_444  =>   energy_bin_pos_data(443 ),
	   o_Energy_Bin_Pos_445  =>   energy_bin_pos_data(444 ),
	   o_Energy_Bin_Pos_446  =>   energy_bin_pos_data(445 ),
	   o_Energy_Bin_Pos_447  =>   energy_bin_pos_data(446 ),
	   o_Energy_Bin_Pos_448  =>   energy_bin_pos_data(447 ),
	   o_Energy_Bin_Pos_449  =>   energy_bin_pos_data(448 ),
	   o_Energy_Bin_Pos_450  =>   energy_bin_pos_data(449 ),
	   o_Energy_Bin_Pos_451  =>   energy_bin_pos_data(450 ),
	   o_Energy_Bin_Pos_452  =>   energy_bin_pos_data(451 ),
	   o_Energy_Bin_Pos_453  =>   energy_bin_pos_data(452 ),
	   o_Energy_Bin_Pos_454  =>   energy_bin_pos_data(453 ),
	   o_Energy_Bin_Pos_455  =>   energy_bin_pos_data(454 ),
	   o_Energy_Bin_Pos_456  =>   energy_bin_pos_data(455 ),
	   o_Energy_Bin_Pos_457  =>   energy_bin_pos_data(456 ),
	   o_Energy_Bin_Pos_458  =>   energy_bin_pos_data(457 ),
	   o_Energy_Bin_Pos_459  =>   energy_bin_pos_data(458 ),
	   o_Energy_Bin_Pos_460  =>   energy_bin_pos_data(459 ),
	   o_Energy_Bin_Pos_461  =>   energy_bin_pos_data(460 ),
	   o_Energy_Bin_Pos_462  =>   energy_bin_pos_data(461 ),
	   o_Energy_Bin_Pos_463  =>   energy_bin_pos_data(462 ),
	   o_Energy_Bin_Pos_464  =>   energy_bin_pos_data(463 ),
	   o_Energy_Bin_Pos_465  =>   energy_bin_pos_data(464 ),
	   o_Energy_Bin_Pos_466  =>   energy_bin_pos_data(465 ),
	   o_Energy_Bin_Pos_467  =>   energy_bin_pos_data(466 ),
	   o_Energy_Bin_Pos_468  =>   energy_bin_pos_data(467 ),
	   o_Energy_Bin_Pos_469  =>   energy_bin_pos_data(468 ),
	   o_Energy_Bin_Pos_470  =>   energy_bin_pos_data(469 ),
	   o_Energy_Bin_Pos_471  =>   energy_bin_pos_data(470 ),
	   o_Energy_Bin_Pos_472  =>   energy_bin_pos_data(471 ),
	   o_Energy_Bin_Pos_473  =>   energy_bin_pos_data(472 ),
	   o_Energy_Bin_Pos_474  =>   energy_bin_pos_data(473 ),
	   o_Energy_Bin_Pos_475  =>   energy_bin_pos_data(474 ),
	   o_Energy_Bin_Pos_476  =>   energy_bin_pos_data(475 ),
	   o_Energy_Bin_Pos_477  =>   energy_bin_pos_data(476 ),
	   o_Energy_Bin_Pos_478  =>   energy_bin_pos_data(477 ),
	   o_Energy_Bin_Pos_479  =>   energy_bin_pos_data(478 ),
	   o_Energy_Bin_Pos_480  =>   energy_bin_pos_data(479 ),
	   o_Energy_Bin_Pos_481  =>   energy_bin_pos_data(480 ),
	   o_Energy_Bin_Pos_482  =>   energy_bin_pos_data(481 ),
	   o_Energy_Bin_Pos_483  =>   energy_bin_pos_data(482 ),
	   o_Energy_Bin_Pos_484  =>   energy_bin_pos_data(483 ),
	   o_Energy_Bin_Pos_485  =>   energy_bin_pos_data(484 ),
	   o_Energy_Bin_Pos_486  =>   energy_bin_pos_data(485 ),
	   o_Energy_Bin_Pos_487  =>   energy_bin_pos_data(486 ),
	   o_Energy_Bin_Pos_488  =>   energy_bin_pos_data(487 ),
	   o_Energy_Bin_Pos_489  =>   energy_bin_pos_data(488 ),
	   o_Energy_Bin_Pos_490  =>   energy_bin_pos_data(489 ),
	   o_Energy_Bin_Pos_491  =>   energy_bin_pos_data(490 ),
	   o_Energy_Bin_Pos_492  =>   energy_bin_pos_data(491 ),
	   o_Energy_Bin_Pos_493  =>   energy_bin_pos_data(492 ),
	   o_Energy_Bin_Pos_494  =>   energy_bin_pos_data(493 ),
	   o_Energy_Bin_Pos_495  =>   energy_bin_pos_data(494 ),
	   o_Energy_Bin_Pos_496  =>   energy_bin_pos_data(495 ),
	   o_Energy_Bin_Pos_497  =>   energy_bin_pos_data(496 ),
	   o_Energy_Bin_Pos_498  =>   energy_bin_pos_data(497 ),
	   o_Energy_Bin_Pos_499  =>   energy_bin_pos_data(498 ),
	   o_Energy_Bin_Pos_500  =>   energy_bin_pos_data(499 ),
	   o_Energy_Bin_Pos_501  =>   energy_bin_pos_data(500 ),
	   o_Energy_Bin_Pos_502  =>   energy_bin_pos_data(501 ),
	   o_Energy_Bin_Pos_503  =>   energy_bin_pos_data(502 ),
	   o_Energy_Bin_Pos_504  =>   energy_bin_pos_data(503 ),
	   o_Energy_Bin_Pos_505  =>   energy_bin_pos_data(504 ),
	   o_Energy_Bin_Pos_506  =>   energy_bin_pos_data(505 ),
	   o_Energy_Bin_Pos_507  =>   energy_bin_pos_data(506 ),
	   o_Energy_Bin_Pos_508  =>   energy_bin_pos_data(507 ),
	   o_Energy_Bin_Pos_509  =>   energy_bin_pos_data(508 ),
	   o_Energy_Bin_Pos_510  =>   energy_bin_pos_data(509 ),
	   o_Energy_Bin_Pos_511  =>   energy_bin_pos_data(510 ),
	   o_Energy_Bin_Pos_512  =>   energy_bin_pos_data(511 ),
	   o_Energy_Bin_Pos_513  =>   energy_bin_pos_data(512 ),
	   o_Energy_Bin_Pos_514  =>   energy_bin_pos_data(513 ),
	   o_Energy_Bin_Pos_515  =>   energy_bin_pos_data(514 ),
	   o_Energy_Bin_Pos_516  =>   energy_bin_pos_data(515 ),
	   o_Energy_Bin_Pos_517  =>   energy_bin_pos_data(516 ),
	   o_Energy_Bin_Pos_518  =>   energy_bin_pos_data(517 ),
	   o_Energy_Bin_Pos_519  =>   energy_bin_pos_data(518 ),
	   o_Energy_Bin_Pos_520  =>   energy_bin_pos_data(519 ),
	   o_Energy_Bin_Pos_521  =>   energy_bin_pos_data(520 ),
	   o_Energy_Bin_Pos_522  =>   energy_bin_pos_data(521 ),
	   o_Energy_Bin_Pos_523  =>   energy_bin_pos_data(522 ),
	   o_Energy_Bin_Pos_524  =>   energy_bin_pos_data(523 ),
	   o_Energy_Bin_Pos_525  =>   energy_bin_pos_data(524 ),
	   o_Energy_Bin_Pos_526  =>   energy_bin_pos_data(525 ),
	   o_Energy_Bin_Pos_527  =>   energy_bin_pos_data(526 ),
	   o_Energy_Bin_Pos_528  =>   energy_bin_pos_data(527 ),
	   o_Energy_Bin_Pos_529  =>   energy_bin_pos_data(528 ),
	   o_Energy_Bin_Pos_530  =>   energy_bin_pos_data(529 ),
	   o_Energy_Bin_Pos_531  =>   energy_bin_pos_data(530 ),
	   o_Energy_Bin_Pos_532  =>   energy_bin_pos_data(531 ),
	   o_Energy_Bin_Pos_533  =>   energy_bin_pos_data(532 ),
	   o_Energy_Bin_Pos_534  =>   energy_bin_pos_data(533 ),
	   o_Energy_Bin_Pos_535  =>   energy_bin_pos_data(534 ),
	   o_Energy_Bin_Pos_536  =>   energy_bin_pos_data(535 ),
	   o_Energy_Bin_Pos_537  =>   energy_bin_pos_data(536 ),
	   o_Energy_Bin_Pos_538  =>   energy_bin_pos_data(537 ),
	   o_Energy_Bin_Pos_539  =>   energy_bin_pos_data(538 ),
	   o_Energy_Bin_Pos_540  =>   energy_bin_pos_data(539 ),
	   o_Energy_Bin_Pos_541  =>   energy_bin_pos_data(540 ),
	   o_Energy_Bin_Pos_542  =>   energy_bin_pos_data(541 ),
	   o_Energy_Bin_Pos_543  =>   energy_bin_pos_data(542 ),
	   o_Energy_Bin_Pos_544  =>   energy_bin_pos_data(543 ),
	   o_Energy_Bin_Pos_545  =>   energy_bin_pos_data(544 ),
	   o_Energy_Bin_Pos_546  =>   energy_bin_pos_data(545 ),
	   o_Energy_Bin_Pos_547  =>   energy_bin_pos_data(546 ),
	   o_Energy_Bin_Pos_548  =>   energy_bin_pos_data(547 ),
	   o_Energy_Bin_Pos_549  =>   energy_bin_pos_data(548 ),
	   o_Energy_Bin_Pos_550  =>   energy_bin_pos_data(549 ),
	   o_Energy_Bin_Pos_551  =>   energy_bin_pos_data(550 ),
	   o_Energy_Bin_Pos_552  =>   energy_bin_pos_data(551 ),
	   o_Energy_Bin_Pos_553  =>   energy_bin_pos_data(552 ),
	   o_Energy_Bin_Pos_554  =>   energy_bin_pos_data(553 ),
	   o_Energy_Bin_Pos_555  =>   energy_bin_pos_data(554 ),
	   o_Energy_Bin_Pos_556  =>   energy_bin_pos_data(555 ),
	   o_Energy_Bin_Pos_557  =>   energy_bin_pos_data(556 ),
	   o_Energy_Bin_Pos_558  =>   energy_bin_pos_data(557 ),
	   o_Energy_Bin_Pos_559  =>   energy_bin_pos_data(558 ),
	   o_Energy_Bin_Pos_560  =>   energy_bin_pos_data(559 ),
	   o_Energy_Bin_Pos_561  =>   energy_bin_pos_data(560 ),
	   o_Energy_Bin_Pos_562  =>   energy_bin_pos_data(561 ),
	   o_Energy_Bin_Pos_563  =>   energy_bin_pos_data(562 ),
	   o_Energy_Bin_Pos_564  =>   energy_bin_pos_data(563 ),
	   o_Energy_Bin_Pos_565  =>   energy_bin_pos_data(564 ),
	   o_Energy_Bin_Pos_566  =>   energy_bin_pos_data(565 ),
	   o_Energy_Bin_Pos_567  =>   energy_bin_pos_data(566 ),
	   o_Energy_Bin_Pos_568  =>   energy_bin_pos_data(567 ),
	   o_Energy_Bin_Pos_569  =>   energy_bin_pos_data(568 ),
	   o_Energy_Bin_Pos_570  =>   energy_bin_pos_data(569 ),
	   o_Energy_Bin_Pos_571  =>   energy_bin_pos_data(570 ),
	   o_Energy_Bin_Pos_572  =>   energy_bin_pos_data(571 ),
	   o_Energy_Bin_Pos_573  =>   energy_bin_pos_data(572 ),
	   o_Energy_Bin_Pos_574  =>   energy_bin_pos_data(573 ),
	   o_Energy_Bin_Pos_575  =>   energy_bin_pos_data(574 ),
	   o_Energy_Bin_Pos_576  =>   energy_bin_pos_data(575 ),
	   o_Energy_Bin_Pos_577  =>   energy_bin_pos_data(576 ),
	   o_Energy_Bin_Pos_578  =>   energy_bin_pos_data(577 ),
	   o_Energy_Bin_Pos_579  =>   energy_bin_pos_data(578 ),
	   o_Energy_Bin_Pos_580  =>   energy_bin_pos_data(579 ),
	   o_Energy_Bin_Pos_581  =>   energy_bin_pos_data(580 ),
	   o_Energy_Bin_Pos_582  =>   energy_bin_pos_data(581 ),
	   o_Energy_Bin_Pos_583  =>   energy_bin_pos_data(582 ),
	   o_Energy_Bin_Pos_584  =>   energy_bin_pos_data(583 ),
	   o_Energy_Bin_Pos_585  =>   energy_bin_pos_data(584 ),
	   o_Energy_Bin_Pos_586  =>   energy_bin_pos_data(585 ),
	   o_Energy_Bin_Pos_587  =>   energy_bin_pos_data(586 ),
	   o_Energy_Bin_Pos_588  =>   energy_bin_pos_data(587 ),
	   o_Energy_Bin_Pos_589  =>   energy_bin_pos_data(588 ),
	   o_Energy_Bin_Pos_590  =>   energy_bin_pos_data(589 ),
	   o_Energy_Bin_Pos_591  =>   energy_bin_pos_data(590 ),
	   o_Energy_Bin_Pos_592  =>   energy_bin_pos_data(591 ),
	   o_Energy_Bin_Pos_593  =>   energy_bin_pos_data(592 ),
	   o_Energy_Bin_Pos_594  =>   energy_bin_pos_data(593 ),
	   o_Energy_Bin_Pos_595  =>   energy_bin_pos_data(594 ),
	   o_Energy_Bin_Pos_596  =>   energy_bin_pos_data(595 ),
	   o_Energy_Bin_Pos_597  =>   energy_bin_pos_data(596 ),
	   o_Energy_Bin_Pos_598  =>   energy_bin_pos_data(597 ),
	   o_Energy_Bin_Pos_599  =>   energy_bin_pos_data(598 ),
	   o_Energy_Bin_Pos_600  =>   energy_bin_pos_data(599 ),
	   o_Energy_Bin_Pos_601  =>   energy_bin_pos_data(600 ),
	   o_Energy_Bin_Pos_602  =>   energy_bin_pos_data(601 ),
	   o_Energy_Bin_Pos_603  =>   energy_bin_pos_data(602 ),
	   o_Energy_Bin_Pos_604  =>   energy_bin_pos_data(603 ),
	   o_Energy_Bin_Pos_605  =>   energy_bin_pos_data(604 ),
	   o_Energy_Bin_Pos_606  =>   energy_bin_pos_data(605 ),
	   o_Energy_Bin_Pos_607  =>   energy_bin_pos_data(606 ),
	   o_Energy_Bin_Pos_608  =>   energy_bin_pos_data(607 ),
	   o_Energy_Bin_Pos_609  =>   energy_bin_pos_data(608 ),
	   o_Energy_Bin_Pos_610  =>   energy_bin_pos_data(609 ),
	   o_Energy_Bin_Pos_611  =>   energy_bin_pos_data(610 ),
	   o_Energy_Bin_Pos_612  =>   energy_bin_pos_data(611 ),
	   o_Energy_Bin_Pos_613  =>   energy_bin_pos_data(612 ),
	   o_Energy_Bin_Pos_614  =>   energy_bin_pos_data(613 ),
	   o_Energy_Bin_Pos_615  =>   energy_bin_pos_data(614 ),
	   o_Energy_Bin_Pos_616  =>   energy_bin_pos_data(615 ),
	   o_Energy_Bin_Pos_617  =>   energy_bin_pos_data(616 ),
	   o_Energy_Bin_Pos_618  =>   energy_bin_pos_data(617 ),
	   o_Energy_Bin_Pos_619  =>   energy_bin_pos_data(618 ),
	   o_Energy_Bin_Pos_620  =>   energy_bin_pos_data(619 ),
	   o_Energy_Bin_Pos_621  =>   energy_bin_pos_data(620 ),
	   o_Energy_Bin_Pos_622  =>   energy_bin_pos_data(621 ),
	   o_Energy_Bin_Pos_623  =>   energy_bin_pos_data(622 ),
	   o_Energy_Bin_Pos_624  =>   energy_bin_pos_data(623 ),
	   o_Energy_Bin_Pos_625  =>   energy_bin_pos_data(624 ),
	   o_Energy_Bin_Pos_626  =>   energy_bin_pos_data(625 ),
	   o_Energy_Bin_Pos_627  =>   energy_bin_pos_data(626 ),
	   o_Energy_Bin_Pos_628  =>   energy_bin_pos_data(627 ),
	   o_Energy_Bin_Pos_629  =>   energy_bin_pos_data(628 ),
	   o_Energy_Bin_Pos_630  =>   energy_bin_pos_data(629 ),
	   o_Energy_Bin_Pos_631  =>   energy_bin_pos_data(630 ),
	   o_Energy_Bin_Pos_632  =>   energy_bin_pos_data(631 ),
	   o_Energy_Bin_Pos_633  =>   energy_bin_pos_data(632 ),
	   o_Energy_Bin_Pos_634  =>   energy_bin_pos_data(633 ),
	   o_Energy_Bin_Pos_635  =>   energy_bin_pos_data(634 ),
	   o_Energy_Bin_Pos_636  =>   energy_bin_pos_data(635 ),
	   o_Energy_Bin_Pos_637  =>   energy_bin_pos_data(636 ),
	   o_Energy_Bin_Pos_638  =>   energy_bin_pos_data(637 ),
	   o_Energy_Bin_Pos_639  =>   energy_bin_pos_data(638 ),
	   o_Energy_Bin_Pos_640  =>   energy_bin_pos_data(639 ),
	   o_Energy_Bin_Pos_641  =>   energy_bin_pos_data(640 ),
	   o_Energy_Bin_Pos_642  =>   energy_bin_pos_data(641 ),
	   o_Energy_Bin_Pos_643  =>   energy_bin_pos_data(642 ),
	   o_Energy_Bin_Pos_644  =>   energy_bin_pos_data(643 ),
	   o_Energy_Bin_Pos_645  =>   energy_bin_pos_data(644 ),
	   o_Energy_Bin_Pos_646  =>   energy_bin_pos_data(645 ),
	   o_Energy_Bin_Pos_647  =>   energy_bin_pos_data(646 ),
	   o_Energy_Bin_Pos_648  =>   energy_bin_pos_data(647 ),
	   o_Energy_Bin_Pos_649  =>   energy_bin_pos_data(648 ),
	   o_Energy_Bin_Pos_650  =>   energy_bin_pos_data(649 ),
	   o_Energy_Bin_Pos_651  =>   energy_bin_pos_data(650 ),
	   o_Energy_Bin_Pos_652  =>   energy_bin_pos_data(651 ),
	   o_Energy_Bin_Pos_653  =>   energy_bin_pos_data(652 ),
	   o_Energy_Bin_Pos_654  =>   energy_bin_pos_data(653 ),
	   o_Energy_Bin_Pos_655  =>   energy_bin_pos_data(654 ),
	   o_Energy_Bin_Pos_656  =>   energy_bin_pos_data(655 ),
	   o_Energy_Bin_Pos_657  =>   energy_bin_pos_data(656 ),
	   o_Energy_Bin_Pos_658  =>   energy_bin_pos_data(657 ),
	   o_Energy_Bin_Pos_659  =>   energy_bin_pos_data(658 ),
	   o_Energy_Bin_Pos_660  =>   energy_bin_pos_data(659 ),
	   o_Energy_Bin_Pos_661  =>   energy_bin_pos_data(660 ),
	   o_Energy_Bin_Pos_662  =>   energy_bin_pos_data(661 ),
	   o_Energy_Bin_Pos_663  =>   energy_bin_pos_data(662 ),
	   o_Energy_Bin_Pos_664  =>   energy_bin_pos_data(663 ),
	   o_Energy_Bin_Pos_665  =>   energy_bin_pos_data(664 ),
	   o_Energy_Bin_Pos_666  =>   energy_bin_pos_data(665 ),
	   o_Energy_Bin_Pos_667  =>   energy_bin_pos_data(666 ),
	   o_Energy_Bin_Pos_668  =>   energy_bin_pos_data(667 ),
	   o_Energy_Bin_Pos_669  =>   energy_bin_pos_data(668 ),
	   o_Energy_Bin_Pos_670  =>   energy_bin_pos_data(669 ),
	   o_Energy_Bin_Pos_671  =>   energy_bin_pos_data(670 ),
	   o_Energy_Bin_Pos_672  =>   energy_bin_pos_data(671 ),
	   o_Energy_Bin_Pos_673  =>   energy_bin_pos_data(672 ),
	   o_Energy_Bin_Pos_674  =>   energy_bin_pos_data(673 ),
	   o_Energy_Bin_Pos_675  =>   energy_bin_pos_data(674 ),
	   o_Energy_Bin_Pos_676  =>   energy_bin_pos_data(675 ),
	   o_Energy_Bin_Pos_677  =>   energy_bin_pos_data(676 ),
	   o_Energy_Bin_Pos_678  =>   energy_bin_pos_data(677 ),
	   o_Energy_Bin_Pos_679  =>   energy_bin_pos_data(678 ),
	   o_Energy_Bin_Pos_680  =>   energy_bin_pos_data(679 ),
	   o_Energy_Bin_Pos_681  =>   energy_bin_pos_data(680 ),
	   o_Energy_Bin_Pos_682  =>   energy_bin_pos_data(681 ),
	   o_Energy_Bin_Pos_683  =>   energy_bin_pos_data(682 ),
	   o_Energy_Bin_Pos_684  =>   energy_bin_pos_data(683 ),
	   o_Energy_Bin_Pos_685  =>   energy_bin_pos_data(684 ),
	   o_Energy_Bin_Pos_686  =>   energy_bin_pos_data(685 ),
	   o_Energy_Bin_Pos_687  =>   energy_bin_pos_data(686 ),
	   o_Energy_Bin_Pos_688  =>   energy_bin_pos_data(687 ),
	   o_Energy_Bin_Pos_689  =>   energy_bin_pos_data(688 ),
	   o_Energy_Bin_Pos_690  =>   energy_bin_pos_data(689 ),
	   o_Energy_Bin_Pos_691  =>   energy_bin_pos_data(690 ),
	   o_Energy_Bin_Pos_692  =>   energy_bin_pos_data(691 ),
	   o_Energy_Bin_Pos_693  =>   energy_bin_pos_data(692 ),
	   o_Energy_Bin_Pos_694  =>   energy_bin_pos_data(693 ),
	   o_Energy_Bin_Pos_695  =>   energy_bin_pos_data(694 ),
	   o_Energy_Bin_Pos_696  =>   energy_bin_pos_data(695 ),
	   o_Energy_Bin_Pos_697  =>   energy_bin_pos_data(696 ),
	   o_Energy_Bin_Pos_698  =>   energy_bin_pos_data(697 ),
	   o_Energy_Bin_Pos_699  =>   energy_bin_pos_data(698 ),
	   o_Energy_Bin_Pos_700  =>   energy_bin_pos_data(699 ),
	   o_Energy_Bin_Pos_701  =>   energy_bin_pos_data(700 ),
	   o_Energy_Bin_Pos_702  =>   energy_bin_pos_data(701 ),
	   o_Energy_Bin_Pos_703  =>   energy_bin_pos_data(702 ),
	   o_Energy_Bin_Pos_704  =>   energy_bin_pos_data(703 ),
	   o_Energy_Bin_Pos_705  =>   energy_bin_pos_data(704 ),
	   o_Energy_Bin_Pos_706  =>   energy_bin_pos_data(705 ),
	   o_Energy_Bin_Pos_707  =>   energy_bin_pos_data(706 ),
	   o_Energy_Bin_Pos_708  =>   energy_bin_pos_data(707 ),
	   o_Energy_Bin_Pos_709  =>   energy_bin_pos_data(708 ),
	   o_Energy_Bin_Pos_710  =>   energy_bin_pos_data(709 ),
	   o_Energy_Bin_Pos_711  =>   energy_bin_pos_data(710 ),
	   o_Energy_Bin_Pos_712  =>   energy_bin_pos_data(711 ),
	   o_Energy_Bin_Pos_713  =>   energy_bin_pos_data(712 ),
	   o_Energy_Bin_Pos_714  =>   energy_bin_pos_data(713 ),
	   o_Energy_Bin_Pos_715  =>   energy_bin_pos_data(714 ),
	   o_Energy_Bin_Pos_716  =>   energy_bin_pos_data(715 ),
	   o_Energy_Bin_Pos_717  =>   energy_bin_pos_data(716 ),
	   o_Energy_Bin_Pos_718  =>   energy_bin_pos_data(717 ),
	   o_Energy_Bin_Pos_719  =>   energy_bin_pos_data(718 ),
	   o_Energy_Bin_Pos_720  =>   energy_bin_pos_data(719 ),
	   o_Energy_Bin_Pos_721  =>   energy_bin_pos_data(720 ),
	   o_Energy_Bin_Pos_722  =>   energy_bin_pos_data(721 ),
	   o_Energy_Bin_Pos_723  =>   energy_bin_pos_data(722 ),
	   o_Energy_Bin_Pos_724  =>   energy_bin_pos_data(723 ),
	   o_Energy_Bin_Pos_725  =>   energy_bin_pos_data(724 ),
	   o_Energy_Bin_Pos_726  =>   energy_bin_pos_data(725 ),
	   o_Energy_Bin_Pos_727  =>   energy_bin_pos_data(726 ),
	   o_Energy_Bin_Pos_728  =>   energy_bin_pos_data(727 ),
	   o_Energy_Bin_Pos_729  =>   energy_bin_pos_data(728 ),
	   o_Energy_Bin_Pos_730  =>   energy_bin_pos_data(729 ),
	   o_Energy_Bin_Pos_731  =>   energy_bin_pos_data(730 ),
	   o_Energy_Bin_Pos_732  =>   energy_bin_pos_data(731 ),
	   o_Energy_Bin_Pos_733  =>   energy_bin_pos_data(732 ),
	   o_Energy_Bin_Pos_734  =>   energy_bin_pos_data(733 ),
	   o_Energy_Bin_Pos_735  =>   energy_bin_pos_data(734 ),
	   o_Energy_Bin_Pos_736  =>   energy_bin_pos_data(735 ),
	   o_Energy_Bin_Pos_737  =>   energy_bin_pos_data(736 ),
	   o_Energy_Bin_Pos_738  =>   energy_bin_pos_data(737 ),
	   o_Energy_Bin_Pos_739  =>   energy_bin_pos_data(738 ),
	   o_Energy_Bin_Pos_740  =>   energy_bin_pos_data(739 ),
	   o_Energy_Bin_Pos_741  =>   energy_bin_pos_data(740 ),
	   o_Energy_Bin_Pos_742  =>   energy_bin_pos_data(741 ),
	   o_Energy_Bin_Pos_743  =>   energy_bin_pos_data(742 ),
	   o_Energy_Bin_Pos_744  =>   energy_bin_pos_data(743 ),
	   o_Energy_Bin_Pos_745  =>   energy_bin_pos_data(744 ),
	   o_Energy_Bin_Pos_746  =>   energy_bin_pos_data(745 ),
	   o_Energy_Bin_Pos_747  =>   energy_bin_pos_data(746 ),
	   o_Energy_Bin_Pos_748  =>   energy_bin_pos_data(747 ),
	   o_Energy_Bin_Pos_749  =>   energy_bin_pos_data(748 ),
	   o_Energy_Bin_Pos_750  =>   energy_bin_pos_data(749 ),
	   o_Energy_Bin_Pos_751  =>   energy_bin_pos_data(750 ),
	   o_Energy_Bin_Pos_752  =>   energy_bin_pos_data(751 ),
	   o_Energy_Bin_Pos_753  =>   energy_bin_pos_data(752 ),
	   o_Energy_Bin_Pos_754  =>   energy_bin_pos_data(753 ),
	   o_Energy_Bin_Pos_755  =>   energy_bin_pos_data(754 ),
	   o_Energy_Bin_Pos_756  =>   energy_bin_pos_data(755 ),
	   o_Energy_Bin_Pos_757  =>   energy_bin_pos_data(756 ),
	   o_Energy_Bin_Pos_758  =>   energy_bin_pos_data(757 ),
	   o_Energy_Bin_Pos_759  =>   energy_bin_pos_data(758 ),
	   o_Energy_Bin_Pos_760  =>   energy_bin_pos_data(759 ),
	   o_Energy_Bin_Pos_761  =>   energy_bin_pos_data(760 ),
	   o_Energy_Bin_Pos_762  =>   energy_bin_pos_data(761 ),
	   o_Energy_Bin_Pos_763  =>   energy_bin_pos_data(762 ),
	   o_Energy_Bin_Pos_764  =>   energy_bin_pos_data(763 ),
	   o_Energy_Bin_Pos_765  =>   energy_bin_pos_data(764 ),
	   o_Energy_Bin_Pos_766  =>   energy_bin_pos_data(765 ),
	   o_Energy_Bin_Pos_767  =>   energy_bin_pos_data(766 ),
	   o_Energy_Bin_Pos_768  =>   energy_bin_pos_data(767 ),
	   o_Energy_Bin_Pos_769  =>   energy_bin_pos_data(768 ),
	   o_Energy_Bin_Pos_770  =>   energy_bin_pos_data(769 ),
	   o_Energy_Bin_Pos_771  =>   energy_bin_pos_data(770 ),
	   o_Energy_Bin_Pos_772  =>   energy_bin_pos_data(771 ),
	   o_Energy_Bin_Pos_773  =>   energy_bin_pos_data(772 ),
	   o_Energy_Bin_Pos_774  =>   energy_bin_pos_data(773 ),
	   o_Energy_Bin_Pos_775  =>   energy_bin_pos_data(774 ),
	   o_Energy_Bin_Pos_776  =>   energy_bin_pos_data(775 ),
	   o_Energy_Bin_Pos_777  =>   energy_bin_pos_data(776 ),
	   o_Energy_Bin_Pos_778  =>   energy_bin_pos_data(777 ),
	   o_Energy_Bin_Pos_779  =>   energy_bin_pos_data(778 ),
	   o_Energy_Bin_Pos_780  =>   energy_bin_pos_data(779 ),
	   o_Energy_Bin_Pos_781  =>   energy_bin_pos_data(780 ),
	   o_Energy_Bin_Pos_782  =>   energy_bin_pos_data(781 ),
	   o_Energy_Bin_Pos_783  =>   energy_bin_pos_data(782 ),
	   o_Energy_Bin_Pos_784  =>   energy_bin_pos_data(783 ),
	   o_Energy_Bin_Pos_785  =>   energy_bin_pos_data(784 ),
	   o_Energy_Bin_Pos_786  =>   energy_bin_pos_data(785 ),
	   o_Energy_Bin_Pos_787  =>   energy_bin_pos_data(786 ),
	   o_Energy_Bin_Pos_788  =>   energy_bin_pos_data(787 ),
	   o_Energy_Bin_Pos_789  =>   energy_bin_pos_data(788 ),
	   o_Energy_Bin_Pos_790  =>   energy_bin_pos_data(789 ),
	   o_Energy_Bin_Pos_791  =>   energy_bin_pos_data(790 ),
	   o_Energy_Bin_Pos_792  =>   energy_bin_pos_data(791 ),
	   o_Energy_Bin_Pos_793  =>   energy_bin_pos_data(792 ),
	   o_Energy_Bin_Pos_794  =>   energy_bin_pos_data(793 ),
	   o_Energy_Bin_Pos_795  =>   energy_bin_pos_data(794 ),
	   o_Energy_Bin_Pos_796  =>   energy_bin_pos_data(795 ),
	   o_Energy_Bin_Pos_797  =>   energy_bin_pos_data(796 ),
	   o_Energy_Bin_Pos_798  =>   energy_bin_pos_data(797 ),
	   o_Energy_Bin_Pos_799  =>   energy_bin_pos_data(798 ),
	   o_Energy_Bin_Pos_800  =>   energy_bin_pos_data(799 ),
	   o_Energy_Bin_Pos_801  =>   energy_bin_pos_data(800 ),
	   o_Energy_Bin_Pos_802  =>   energy_bin_pos_data(801 ),
	   o_Energy_Bin_Pos_803  =>   energy_bin_pos_data(802 ),
	   o_Energy_Bin_Pos_804  =>   energy_bin_pos_data(803 ),
	   o_Energy_Bin_Pos_805  =>   energy_bin_pos_data(804 ),
	   o_Energy_Bin_Pos_806  =>   energy_bin_pos_data(805 ),
	   o_Energy_Bin_Pos_807  =>   energy_bin_pos_data(806 ),
	   o_Energy_Bin_Pos_808  =>   energy_bin_pos_data(807 ),
	   o_Energy_Bin_Pos_809  =>   energy_bin_pos_data(808 ),
	   o_Energy_Bin_Pos_810  =>   energy_bin_pos_data(809 ),
	   o_Energy_Bin_Pos_811  =>   energy_bin_pos_data(810 ),
	   o_Energy_Bin_Pos_812  =>   energy_bin_pos_data(811 ),
	   o_Energy_Bin_Pos_813  =>   energy_bin_pos_data(812 ),
	   o_Energy_Bin_Pos_814  =>   energy_bin_pos_data(813 ),
	   o_Energy_Bin_Pos_815  =>   energy_bin_pos_data(814 ),
	   o_Energy_Bin_Pos_816  =>   energy_bin_pos_data(815 ),
	   o_Energy_Bin_Pos_817  =>   energy_bin_pos_data(816 ),
	   o_Energy_Bin_Pos_818  =>   energy_bin_pos_data(817 ),
	   o_Energy_Bin_Pos_819  =>   energy_bin_pos_data(818 ),
	   o_Energy_Bin_Pos_820  =>   energy_bin_pos_data(819 ),
	   o_Energy_Bin_Pos_821  =>   energy_bin_pos_data(820 ),
	   o_Energy_Bin_Pos_822  =>   energy_bin_pos_data(821 ),
	   o_Energy_Bin_Pos_823  =>   energy_bin_pos_data(822 ),
	   o_Energy_Bin_Pos_824  =>   energy_bin_pos_data(823 ),
	   o_Energy_Bin_Pos_825  =>   energy_bin_pos_data(824 ),
	   o_Energy_Bin_Pos_826  =>   energy_bin_pos_data(825 ),
	   o_Energy_Bin_Pos_827  =>   energy_bin_pos_data(826 ),
	   o_Energy_Bin_Pos_828  =>   energy_bin_pos_data(827 ),
	   o_Energy_Bin_Pos_829  =>   energy_bin_pos_data(828 ),
	   o_Energy_Bin_Pos_830  =>   energy_bin_pos_data(829 ),
	   o_Energy_Bin_Pos_831  =>   energy_bin_pos_data(830 ),
	   o_Energy_Bin_Pos_832  =>   energy_bin_pos_data(831 ),
	   o_Energy_Bin_Pos_833  =>   energy_bin_pos_data(832 ),
	   o_Energy_Bin_Pos_834  =>   energy_bin_pos_data(833 ),
	   o_Energy_Bin_Pos_835  =>   energy_bin_pos_data(834 ),
	   o_Energy_Bin_Pos_836  =>   energy_bin_pos_data(835 ),
	   o_Energy_Bin_Pos_837  =>   energy_bin_pos_data(836 ),
	   o_Energy_Bin_Pos_838  =>   energy_bin_pos_data(837 ),
	   o_Energy_Bin_Pos_839  =>   energy_bin_pos_data(838 ),
	   o_Energy_Bin_Pos_840  =>   energy_bin_pos_data(839 ),
	   o_Energy_Bin_Pos_841  =>   energy_bin_pos_data(840 ),
	   o_Energy_Bin_Pos_842  =>   energy_bin_pos_data(841 ),
	   o_Energy_Bin_Pos_843  =>   energy_bin_pos_data(842 ),
	   o_Energy_Bin_Pos_844  =>   energy_bin_pos_data(843 ),
	   o_Energy_Bin_Pos_845  =>   energy_bin_pos_data(844 ),
	   o_Energy_Bin_Pos_846  =>   energy_bin_pos_data(845 ),
	   o_Energy_Bin_Pos_847  =>   energy_bin_pos_data(846 ),
	   o_Energy_Bin_Pos_848  =>   energy_bin_pos_data(847 ),
	   o_Energy_Bin_Pos_849  =>   energy_bin_pos_data(848 ),
	   o_Energy_Bin_Pos_850  =>   energy_bin_pos_data(849 ),
	   o_Energy_Bin_Pos_851  =>   energy_bin_pos_data(850 ),
	   o_Energy_Bin_Pos_852  =>   energy_bin_pos_data(851 ),
	   o_Energy_Bin_Pos_853  =>   energy_bin_pos_data(852 ),
	   o_Energy_Bin_Pos_854  =>   energy_bin_pos_data(853 ),
	   o_Energy_Bin_Pos_855  =>   energy_bin_pos_data(854 ),
	   o_Energy_Bin_Pos_856  =>   energy_bin_pos_data(855 ),
	   o_Energy_Bin_Pos_857  =>   energy_bin_pos_data(856 ),
	   o_Energy_Bin_Pos_858  =>   energy_bin_pos_data(857 ),
	   o_Energy_Bin_Pos_859  =>   energy_bin_pos_data(858 ),
	   o_Energy_Bin_Pos_860  =>   energy_bin_pos_data(859 ),
	   o_Energy_Bin_Pos_861  =>   energy_bin_pos_data(860 ),
	   o_Energy_Bin_Pos_862  =>   energy_bin_pos_data(861 ),
	   o_Energy_Bin_Pos_863  =>   energy_bin_pos_data(862 ),
	   o_Energy_Bin_Pos_864  =>   energy_bin_pos_data(863 ),
	   o_Energy_Bin_Pos_865  =>   energy_bin_pos_data(864 ),
	   o_Energy_Bin_Pos_866  =>   energy_bin_pos_data(865 ),
	   o_Energy_Bin_Pos_867  =>   energy_bin_pos_data(866 ),
	   o_Energy_Bin_Pos_868  =>   energy_bin_pos_data(867 ),
	   o_Energy_Bin_Pos_869  =>   energy_bin_pos_data(868 ),
	   o_Energy_Bin_Pos_870  =>   energy_bin_pos_data(869 ),
	   o_Energy_Bin_Pos_871  =>   energy_bin_pos_data(870 ),
	   o_Energy_Bin_Pos_872  =>   energy_bin_pos_data(871 ),
	   o_Energy_Bin_Pos_873  =>   energy_bin_pos_data(872 ),
	   o_Energy_Bin_Pos_874  =>   energy_bin_pos_data(873 ),
	   o_Energy_Bin_Pos_875  =>   energy_bin_pos_data(874 ),
	   o_Energy_Bin_Pos_876  =>   energy_bin_pos_data(875 ),
	   o_Energy_Bin_Pos_877  =>   energy_bin_pos_data(876 ),
	   o_Energy_Bin_Pos_878  =>   energy_bin_pos_data(877 ),
	   o_Energy_Bin_Pos_879  =>   energy_bin_pos_data(878 ),
	   o_Energy_Bin_Pos_880  =>   energy_bin_pos_data(879 ),
	   o_Energy_Bin_Pos_881  =>   energy_bin_pos_data(880 ),
	   o_Energy_Bin_Pos_882  =>   energy_bin_pos_data(881 ),
	   o_Energy_Bin_Pos_883  =>   energy_bin_pos_data(882 ),
	   o_Energy_Bin_Pos_884  =>   energy_bin_pos_data(883 ),
	   o_Energy_Bin_Pos_885  =>   energy_bin_pos_data(884 ),
	   o_Energy_Bin_Pos_886  =>   energy_bin_pos_data(885 ),
	   o_Energy_Bin_Pos_887  =>   energy_bin_pos_data(886 ),
	   o_Energy_Bin_Pos_888  =>   energy_bin_pos_data(887 ),
	   o_Energy_Bin_Pos_889  =>   energy_bin_pos_data(888 ),
	   o_Energy_Bin_Pos_890  =>   energy_bin_pos_data(889 ),
	   o_Energy_Bin_Pos_891  =>   energy_bin_pos_data(890 ),
	   o_Energy_Bin_Pos_892  =>   energy_bin_pos_data(891 ),
	   o_Energy_Bin_Pos_893  =>   energy_bin_pos_data(892 ),
	   o_Energy_Bin_Pos_894  =>   energy_bin_pos_data(893 ),
	   o_Energy_Bin_Pos_895  =>   energy_bin_pos_data(894 ),
	   o_Energy_Bin_Pos_896  =>   energy_bin_pos_data(895 ),
	   o_Energy_Bin_Pos_897  =>   energy_bin_pos_data(896 ),
	   o_Energy_Bin_Pos_898  =>   energy_bin_pos_data(897 ),
	   o_Energy_Bin_Pos_899  =>   energy_bin_pos_data(898 ),
	   o_Energy_Bin_Pos_900  =>   energy_bin_pos_data(899 ),
	   o_Energy_Bin_Pos_901  =>   energy_bin_pos_data(900 ),
	   o_Energy_Bin_Pos_902  =>   energy_bin_pos_data(901 ),
	   o_Energy_Bin_Pos_903  =>   energy_bin_pos_data(902 ),
	   o_Energy_Bin_Pos_904  =>   energy_bin_pos_data(903 ),
	   o_Energy_Bin_Pos_905  =>   energy_bin_pos_data(904 ),
	   o_Energy_Bin_Pos_906  =>   energy_bin_pos_data(905 ),
	   o_Energy_Bin_Pos_907  =>   energy_bin_pos_data(906 ),
	   o_Energy_Bin_Pos_908  =>   energy_bin_pos_data(907 ),
	   o_Energy_Bin_Pos_909  =>   energy_bin_pos_data(908 ),
	   o_Energy_Bin_Pos_910  =>   energy_bin_pos_data(909 ),
	   o_Energy_Bin_Pos_911  =>   energy_bin_pos_data(910 ),
	   o_Energy_Bin_Pos_912  =>   energy_bin_pos_data(911 ),
	   o_Energy_Bin_Pos_913  =>   energy_bin_pos_data(912 ),
	   o_Energy_Bin_Pos_914  =>   energy_bin_pos_data(913 ),
	   o_Energy_Bin_Pos_915  =>   energy_bin_pos_data(914 ),
	   o_Energy_Bin_Pos_916  =>   energy_bin_pos_data(915 ),
	   o_Energy_Bin_Pos_917  =>   energy_bin_pos_data(916 ),
	   o_Energy_Bin_Pos_918  =>   energy_bin_pos_data(917 ),
	   o_Energy_Bin_Pos_919  =>   energy_bin_pos_data(918 ),
	   o_Energy_Bin_Pos_920  =>   energy_bin_pos_data(919 ),
	   o_Energy_Bin_Pos_921  =>   energy_bin_pos_data(920 ),
	   o_Energy_Bin_Pos_922  =>   energy_bin_pos_data(921 ),
	   o_Energy_Bin_Pos_923  =>   energy_bin_pos_data(922 ),
	   o_Energy_Bin_Pos_924  =>   energy_bin_pos_data(923 ),
	   o_Energy_Bin_Pos_925  =>   energy_bin_pos_data(924 ),
	   o_Energy_Bin_Pos_926  =>   energy_bin_pos_data(925 ),
	   o_Energy_Bin_Pos_927  =>   energy_bin_pos_data(926 ),
	   o_Energy_Bin_Pos_928  =>   energy_bin_pos_data(927 ),
	   o_Energy_Bin_Pos_929  =>   energy_bin_pos_data(928 ),
	   o_Energy_Bin_Pos_930  =>   energy_bin_pos_data(929 ),
	   o_Energy_Bin_Pos_931  =>   energy_bin_pos_data(930 ),
	   o_Energy_Bin_Pos_932  =>   energy_bin_pos_data(931 ),
	   o_Energy_Bin_Pos_933  =>   energy_bin_pos_data(932 ),
	   o_Energy_Bin_Pos_934  =>   energy_bin_pos_data(933 ),
	   o_Energy_Bin_Pos_935  =>   energy_bin_pos_data(934 ),
	   o_Energy_Bin_Pos_936  =>   energy_bin_pos_data(935 ),
	   o_Energy_Bin_Pos_937  =>   energy_bin_pos_data(936 ),
	   o_Energy_Bin_Pos_938  =>   energy_bin_pos_data(937 ),
	   o_Energy_Bin_Pos_939  =>   energy_bin_pos_data(938 ),
	   o_Energy_Bin_Pos_940  =>   energy_bin_pos_data(939 ),
	   o_Energy_Bin_Pos_941  =>   energy_bin_pos_data(940 ),
	   o_Energy_Bin_Pos_942  =>   energy_bin_pos_data(941 ),
	   o_Energy_Bin_Pos_943  =>   energy_bin_pos_data(942 ),
	   o_Energy_Bin_Pos_944  =>   energy_bin_pos_data(943 ),
	   o_Energy_Bin_Pos_945  =>   energy_bin_pos_data(944 ),
	   o_Energy_Bin_Pos_946  =>   energy_bin_pos_data(945 ),
	   o_Energy_Bin_Pos_947  =>   energy_bin_pos_data(946 ),
	   o_Energy_Bin_Pos_948  =>   energy_bin_pos_data(947 ),
	   o_Energy_Bin_Pos_949  =>   energy_bin_pos_data(948 ),
	   o_Energy_Bin_Pos_950  =>   energy_bin_pos_data(949 ),
	   o_Energy_Bin_Pos_951  =>   energy_bin_pos_data(950 ),
	   o_Energy_Bin_Pos_952  =>   energy_bin_pos_data(951 ),
	   o_Energy_Bin_Pos_953  =>   energy_bin_pos_data(952 ),
	   o_Energy_Bin_Pos_954  =>   energy_bin_pos_data(953 ),
	   o_Energy_Bin_Pos_955  =>   energy_bin_pos_data(954 ),
	   o_Energy_Bin_Pos_956  =>   energy_bin_pos_data(955 ),
	   o_Energy_Bin_Pos_957  =>   energy_bin_pos_data(956 ),
	   o_Energy_Bin_Pos_958  =>   energy_bin_pos_data(957 ),
	   o_Energy_Bin_Pos_959  =>   energy_bin_pos_data(958 ),
	   o_Energy_Bin_Pos_960  =>   energy_bin_pos_data(959 ),
	   o_Energy_Bin_Pos_961  =>   energy_bin_pos_data(960 ),
	   o_Energy_Bin_Pos_962  =>   energy_bin_pos_data(961 ),
	   o_Energy_Bin_Pos_963  =>   energy_bin_pos_data(962 ),
	   o_Energy_Bin_Pos_964  =>   energy_bin_pos_data(963 ),
	   o_Energy_Bin_Pos_965  =>   energy_bin_pos_data(964 ),
	   o_Energy_Bin_Pos_966  =>   energy_bin_pos_data(965 ),
	   o_Energy_Bin_Pos_967  =>   energy_bin_pos_data(966 ),
	   o_Energy_Bin_Pos_968  =>   energy_bin_pos_data(967 ),
	   o_Energy_Bin_Pos_969  =>   energy_bin_pos_data(968 ),
	   o_Energy_Bin_Pos_970  =>   energy_bin_pos_data(969 ),
	   o_Energy_Bin_Pos_971  =>   energy_bin_pos_data(970 ),
	   o_Energy_Bin_Pos_972  =>   energy_bin_pos_data(971 ),
	   o_Energy_Bin_Pos_973  =>   energy_bin_pos_data(972 ),
	   o_Energy_Bin_Pos_974  =>   energy_bin_pos_data(973 ),
	   o_Energy_Bin_Pos_975  =>   energy_bin_pos_data(974 ),
	   o_Energy_Bin_Pos_976  =>   energy_bin_pos_data(975 ),
	   o_Energy_Bin_Pos_977  =>   energy_bin_pos_data(976 ),
	   o_Energy_Bin_Pos_978  =>   energy_bin_pos_data(977 ),
	   o_Energy_Bin_Pos_979  =>   energy_bin_pos_data(978 ),
	   o_Energy_Bin_Pos_980  =>   energy_bin_pos_data(979 ),
	   o_Energy_Bin_Pos_981  =>   energy_bin_pos_data(980 ),
	   o_Energy_Bin_Pos_982  =>   energy_bin_pos_data(981 ),
	   o_Energy_Bin_Pos_983  =>   energy_bin_pos_data(982 ),
	   o_Energy_Bin_Pos_984  =>   energy_bin_pos_data(983 ),
	   o_Energy_Bin_Pos_985  =>   energy_bin_pos_data(984 ),
	   o_Energy_Bin_Pos_986  =>   energy_bin_pos_data(985 ),
	   o_Energy_Bin_Pos_987  =>   energy_bin_pos_data(986 ),
	   o_Energy_Bin_Pos_988  =>   energy_bin_pos_data(987 ),
	   o_Energy_Bin_Pos_989  =>   energy_bin_pos_data(988 ),
	   o_Energy_Bin_Pos_990  =>   energy_bin_pos_data(989 ),
	   o_Energy_Bin_Pos_991  =>   energy_bin_pos_data(990 ),
	   o_Energy_Bin_Pos_992  =>   energy_bin_pos_data(991 ),
	   o_Energy_Bin_Pos_993  =>   energy_bin_pos_data(992 ),
	   o_Energy_Bin_Pos_994  =>   energy_bin_pos_data(993 ),
	   o_Energy_Bin_Pos_995  =>   energy_bin_pos_data(994 ),
	   o_Energy_Bin_Pos_996  =>   energy_bin_pos_data(995 ),
	   o_Energy_Bin_Pos_997  =>   energy_bin_pos_data(996 ),
	   o_Energy_Bin_Pos_998  =>   energy_bin_pos_data(997 ),
	   o_Energy_Bin_Pos_999  =>   energy_bin_pos_data(998 ),
	   o_Energy_Bin_Pos_1000 =>   energy_bin_pos_data(999 ),
	   o_Energy_Bin_Pos_1001 =>   energy_bin_pos_data(1000),
	   o_Energy_Bin_Pos_1002 =>   energy_bin_pos_data(1001),
	   o_Energy_Bin_Pos_1003 =>   energy_bin_pos_data(1002),
	   o_Energy_Bin_Pos_1004 =>   energy_bin_pos_data(1003),
	   o_Energy_Bin_Pos_1005 =>   energy_bin_pos_data(1004),
	   o_Energy_Bin_Pos_1006 =>   energy_bin_pos_data(1005),
	   o_Energy_Bin_Pos_1007 =>   energy_bin_pos_data(1006),
	   o_Energy_Bin_Pos_1008 =>   energy_bin_pos_data(1007),
	   o_Energy_Bin_Pos_1009 =>   energy_bin_pos_data(1008),
	   o_Energy_Bin_Pos_1010 =>   energy_bin_pos_data(1009),
	   o_Energy_Bin_Pos_1011 =>   energy_bin_pos_data(1010),
	   o_Energy_Bin_Pos_1012 =>   energy_bin_pos_data(1011),
	   o_Energy_Bin_Pos_1013 =>   energy_bin_pos_data(1012),
	   o_Energy_Bin_Pos_1014 =>   energy_bin_pos_data(1013),
	   o_Energy_Bin_Pos_1015 =>   energy_bin_pos_data(1014),
	   o_Energy_Bin_Pos_1016 =>   energy_bin_pos_data(1015),
	   o_Energy_Bin_Pos_1017 =>   energy_bin_pos_data(1016),
	   o_Energy_Bin_Pos_1018 =>   energy_bin_pos_data(1017),
	   o_Energy_Bin_Pos_1019 =>   energy_bin_pos_data(1018),
	   o_Energy_Bin_Pos_1020 =>   energy_bin_pos_data(1019),
	   o_Energy_Bin_Pos_1021 =>   energy_bin_pos_data(1020),
	   o_Energy_Bin_Pos_1022 =>   energy_bin_pos_data(1021),
	   o_Energy_Bin_Pos_1023 =>   energy_bin_pos_data(1022),
	   o_Energy_Bin_Pos_1024 =>   energy_bin_pos_data(1023),	   
	   
	   o_Energy_Bin_1        =>   energy_bin_neg_data(0	  ),
	   o_Energy_Bin_2        =>   energy_bin_neg_data(1   ),
	   o_Energy_Bin_3        =>   energy_bin_neg_data(2   ),
	   o_Energy_Bin_4        =>   energy_bin_neg_data(3   ),
	   o_Energy_Bin_5        =>   energy_bin_neg_data(4   ),
	   o_Energy_Bin_6        =>   energy_bin_neg_data(5   ),
	   o_Energy_Bin_7        =>   energy_bin_neg_data(6   ),
	   o_Energy_Bin_8        =>   energy_bin_neg_data(7   ),
	   o_Energy_Bin_9        =>   energy_bin_neg_data(8   ),
	   o_Energy_Bin_10       =>   energy_bin_neg_data(9   ),
	   o_Energy_Bin_11       =>   energy_bin_neg_data(10  ),
	   o_Energy_Bin_12       =>   energy_bin_neg_data(11  ),
	   o_Energy_Bin_13       =>   energy_bin_neg_data(12  ),
	   o_Energy_Bin_14       =>   energy_bin_neg_data(13  ),
	   o_Energy_Bin_15       =>   energy_bin_neg_data(14  ),
	   o_Energy_Bin_16       =>   energy_bin_neg_data(15  ),
	   o_Energy_Bin_17       =>   energy_bin_neg_data(16  ),
	   o_Energy_Bin_18       =>   energy_bin_neg_data(17  ),
	   o_Energy_Bin_19       =>   energy_bin_neg_data(18  ),
	   o_Energy_Bin_20       =>   energy_bin_neg_data(19  ),
	   o_Energy_Bin_21       =>   energy_bin_neg_data(20  ),
	   o_Energy_Bin_22       =>   energy_bin_neg_data(21  ),
	   o_Energy_Bin_23       =>   energy_bin_neg_data(22  ),
	   o_Energy_Bin_24       =>   energy_bin_neg_data(23  ),
	   o_Energy_Bin_25       =>   energy_bin_neg_data(24  ),
	   o_Energy_Bin_26       =>   energy_bin_neg_data(25  ),
	   o_Energy_Bin_27       =>   energy_bin_neg_data(26  ),
	   o_Energy_Bin_28       =>   energy_bin_neg_data(27  ),
	   o_Energy_Bin_29       =>   energy_bin_neg_data(28  ),
	   o_Energy_Bin_30       =>   energy_bin_neg_data(29  ),
	   o_Energy_Bin_31       =>   energy_bin_neg_data(30  ),
	   o_Energy_Bin_32       =>   energy_bin_neg_data(31  ),
	   o_Energy_Bin_33       =>   energy_bin_neg_data(32  ),
	   o_Energy_Bin_34       =>   energy_bin_neg_data(33  ),
	   o_Energy_Bin_35       =>   energy_bin_neg_data(34  ),
	   o_Energy_Bin_36       =>   energy_bin_neg_data(35  ),
	   o_Energy_Bin_37       =>   energy_bin_neg_data(36  ),
	   o_Energy_Bin_38       =>   energy_bin_neg_data(37  ),
	   o_Energy_Bin_39       =>   energy_bin_neg_data(38  ),
	   o_Energy_Bin_40       =>   energy_bin_neg_data(39  ),
	   o_Energy_Bin_41       =>   energy_bin_neg_data(40  ),
	   o_Energy_Bin_42       =>   energy_bin_neg_data(41  ),
	   o_Energy_Bin_43       =>   energy_bin_neg_data(42  ),
	   o_Energy_Bin_44       =>   energy_bin_neg_data(43  ),
	   o_Energy_Bin_45       =>   energy_bin_neg_data(44  ),
	   o_Energy_Bin_46       =>   energy_bin_neg_data(45  ),
	   o_Energy_Bin_47       =>   energy_bin_neg_data(46  ),
	   o_Energy_Bin_48       =>   energy_bin_neg_data(47  ),
	   o_Energy_Bin_49       =>   energy_bin_neg_data(48  ),
	   o_Energy_Bin_50       =>   energy_bin_neg_data(49  ),
	   o_Energy_Bin_51       =>   energy_bin_neg_data(50  ),
	   o_Energy_Bin_52       =>   energy_bin_neg_data(51  ),
	   o_Energy_Bin_53       =>   energy_bin_neg_data(52  ),
	   o_Energy_Bin_54       =>   energy_bin_neg_data(53  ),
	   o_Energy_Bin_55       =>   energy_bin_neg_data(54  ),
	   o_Energy_Bin_56       =>   energy_bin_neg_data(55  ),
	   o_Energy_Bin_57       =>   energy_bin_neg_data(56  ),
	   o_Energy_Bin_58       =>   energy_bin_neg_data(57  ),
	   o_Energy_Bin_59       =>   energy_bin_neg_data(58  ),
	   o_Energy_Bin_60       =>   energy_bin_neg_data(59  ),
	   o_Energy_Bin_61       =>   energy_bin_neg_data(60  ),
	   o_Energy_Bin_62       =>   energy_bin_neg_data(61  ),
	   o_Energy_Bin_63       =>   energy_bin_neg_data(62  ),
	   o_Energy_Bin_64       =>   energy_bin_neg_data(63  ),
	   o_Energy_Bin_65       =>   energy_bin_neg_data(64  ),
	   o_Energy_Bin_66       =>   energy_bin_neg_data(65  ),
	   o_Energy_Bin_67       =>   energy_bin_neg_data(66  ),
	   o_Energy_Bin_68       =>   energy_bin_neg_data(67  ),
	   o_Energy_Bin_69       =>   energy_bin_neg_data(68  ),
	   o_Energy_Bin_70       =>   energy_bin_neg_data(69  ),
	   o_Energy_Bin_71       =>   energy_bin_neg_data(70  ),
	   o_Energy_Bin_72       =>   energy_bin_neg_data(71  ),
	   o_Energy_Bin_73       =>   energy_bin_neg_data(72  ),
	   o_Energy_Bin_74       =>   energy_bin_neg_data(73  ),
	   o_Energy_Bin_75       =>   energy_bin_neg_data(74  ),
	   o_Energy_Bin_76       =>   energy_bin_neg_data(75  ),
	   o_Energy_Bin_77       =>   energy_bin_neg_data(76  ),
	   o_Energy_Bin_78       =>   energy_bin_neg_data(77  ),
	   o_Energy_Bin_79       =>   energy_bin_neg_data(78  ),
	   o_Energy_Bin_80       =>   energy_bin_neg_data(79  ),
	   o_Energy_Bin_81       =>   energy_bin_neg_data(80  ),
	   o_Energy_Bin_82       =>   energy_bin_neg_data(81  ),
	   o_Energy_Bin_83       =>   energy_bin_neg_data(82  ),
	   o_Energy_Bin_84       =>   energy_bin_neg_data(83  ),
	   o_Energy_Bin_85       =>   energy_bin_neg_data(84  ),
	   o_Energy_Bin_86       =>   energy_bin_neg_data(85  ),
	   o_Energy_Bin_87       =>   energy_bin_neg_data(86  ),
	   o_Energy_Bin_88       =>   energy_bin_neg_data(87  ),
	   o_Energy_Bin_89       =>   energy_bin_neg_data(88  ),
	   o_Energy_Bin_90       =>   energy_bin_neg_data(89  ),
	   o_Energy_Bin_91       =>   energy_bin_neg_data(90  ),
	   o_Energy_Bin_92       =>   energy_bin_neg_data(91  ),
	   o_Energy_Bin_93       =>   energy_bin_neg_data(92  ),
	   o_Energy_Bin_94       =>   energy_bin_neg_data(93  ),
	   o_Energy_Bin_95       =>   energy_bin_neg_data(94  ),
	   o_Energy_Bin_96       =>   energy_bin_neg_data(95  ),
	   o_Energy_Bin_97       =>   energy_bin_neg_data(96  ),
	   o_Energy_Bin_98       =>   energy_bin_neg_data(97  ),
	   o_Energy_Bin_99       =>   energy_bin_neg_data(98  ),
	   o_Energy_Bin_100      =>   energy_bin_neg_data(99  ),
	   o_Energy_Bin_101      =>   energy_bin_neg_data(100 ),
	   o_Energy_Bin_102      =>   energy_bin_neg_data(101 ),
	   o_Energy_Bin_103      =>   energy_bin_neg_data(102 ),
	   o_Energy_Bin_104      =>   energy_bin_neg_data(103 ),
	   o_Energy_Bin_105      =>   energy_bin_neg_data(104 ),
	   o_Energy_Bin_106      =>   energy_bin_neg_data(105 ),
	   o_Energy_Bin_107      =>   energy_bin_neg_data(106 ),
	   o_Energy_Bin_108      =>   energy_bin_neg_data(107 ),
	   o_Energy_Bin_109      =>   energy_bin_neg_data(108 ),
	   o_Energy_Bin_110      =>   energy_bin_neg_data(109 ),
	   o_Energy_Bin_111      =>   energy_bin_neg_data(110 ),
	   o_Energy_Bin_112      =>   energy_bin_neg_data(111 ),
	   o_Energy_Bin_113      =>   energy_bin_neg_data(112 ),
	   o_Energy_Bin_114      =>   energy_bin_neg_data(113 ),
	   o_Energy_Bin_115      =>   energy_bin_neg_data(114 ),
	   o_Energy_Bin_116      =>   energy_bin_neg_data(115 ),
	   o_Energy_Bin_117      =>   energy_bin_neg_data(116 ),
	   o_Energy_Bin_118      =>   energy_bin_neg_data(117 ),
	   o_Energy_Bin_119      =>   energy_bin_neg_data(118 ),
	   o_Energy_Bin_120      =>   energy_bin_neg_data(119 ),
	   o_Energy_Bin_121      =>   energy_bin_neg_data(120 ),
	   o_Energy_Bin_122      =>   energy_bin_neg_data(121 ),
	   o_Energy_Bin_123      =>   energy_bin_neg_data(122 ),
	   o_Energy_Bin_124      =>   energy_bin_neg_data(123 ),
	   o_Energy_Bin_125      =>   energy_bin_neg_data(124 ),
	   o_Energy_Bin_126      =>   energy_bin_neg_data(125 ),
	   o_Energy_Bin_127      =>   energy_bin_neg_data(126 ),
	   o_Energy_Bin_128      =>   energy_bin_neg_data(127 ),
	   o_Energy_Bin_129      =>   energy_bin_neg_data(128 ),
	   o_Energy_Bin_130      =>   energy_bin_neg_data(129 ),
	   o_Energy_Bin_131      =>   energy_bin_neg_data(130 ),
	   o_Energy_Bin_132      =>   energy_bin_neg_data(131 ),
	   o_Energy_Bin_133      =>   energy_bin_neg_data(132 ),
	   o_Energy_Bin_134      =>   energy_bin_neg_data(133 ),
	   o_Energy_Bin_135      =>   energy_bin_neg_data(134 ),
	   o_Energy_Bin_136      =>   energy_bin_neg_data(135 ),
	   o_Energy_Bin_137      =>   energy_bin_neg_data(136 ),
	   o_Energy_Bin_138      =>   energy_bin_neg_data(137 ),
	   o_Energy_Bin_139      =>   energy_bin_neg_data(138 ),
	   o_Energy_Bin_140      =>   energy_bin_neg_data(139 ),
	   o_Energy_Bin_141      =>   energy_bin_neg_data(140 ),
	   o_Energy_Bin_142      =>   energy_bin_neg_data(141 ),
	   o_Energy_Bin_143      =>   energy_bin_neg_data(142 ),
	   o_Energy_Bin_144      =>   energy_bin_neg_data(143 ),
	   o_Energy_Bin_145      =>   energy_bin_neg_data(144 ),
	   o_Energy_Bin_146      =>   energy_bin_neg_data(145 ),
	   o_Energy_Bin_147      =>   energy_bin_neg_data(146 ),
	   o_Energy_Bin_148      =>   energy_bin_neg_data(147 ),
	   o_Energy_Bin_149      =>   energy_bin_neg_data(148 ),
	   o_Energy_Bin_150      =>   energy_bin_neg_data(149 ),
	   o_Energy_Bin_151      =>   energy_bin_neg_data(150 ),
	   o_Energy_Bin_152      =>   energy_bin_neg_data(151 ),
	   o_Energy_Bin_153      =>   energy_bin_neg_data(152 ),
	   o_Energy_Bin_154      =>   energy_bin_neg_data(153 ),
	   o_Energy_Bin_155      =>   energy_bin_neg_data(154 ),
	   o_Energy_Bin_156      =>   energy_bin_neg_data(155 ),
	   o_Energy_Bin_157      =>   energy_bin_neg_data(156 ),
	   o_Energy_Bin_158      =>   energy_bin_neg_data(157 ),
	   o_Energy_Bin_159      =>   energy_bin_neg_data(158 ),
	   o_Energy_Bin_160      =>   energy_bin_neg_data(159 ),
	   o_Energy_Bin_161      =>   energy_bin_neg_data(160 ),
	   o_Energy_Bin_162      =>   energy_bin_neg_data(161 ),
	   o_Energy_Bin_163      =>   energy_bin_neg_data(162 ),
	   o_Energy_Bin_164      =>   energy_bin_neg_data(163 ),
	   o_Energy_Bin_165      =>   energy_bin_neg_data(164 ),
	   o_Energy_Bin_166      =>   energy_bin_neg_data(165 ),
	   o_Energy_Bin_167      =>   energy_bin_neg_data(166 ),
	   o_Energy_Bin_168      =>   energy_bin_neg_data(167 ),
	   o_Energy_Bin_169      =>   energy_bin_neg_data(168 ),
	   o_Energy_Bin_170      =>   energy_bin_neg_data(169 ),
	   o_Energy_Bin_171      =>   energy_bin_neg_data(170 ),
	   o_Energy_Bin_172      =>   energy_bin_neg_data(171 ),
	   o_Energy_Bin_173      =>   energy_bin_neg_data(172 ),
	   o_Energy_Bin_174      =>   energy_bin_neg_data(173 ),
	   o_Energy_Bin_175      =>   energy_bin_neg_data(174 ),
	   o_Energy_Bin_176      =>   energy_bin_neg_data(175 ),
	   o_Energy_Bin_177      =>   energy_bin_neg_data(176 ),
	   o_Energy_Bin_178      =>   energy_bin_neg_data(177 ),
	   o_Energy_Bin_179      =>   energy_bin_neg_data(178 ),
	   o_Energy_Bin_180      =>   energy_bin_neg_data(179 ),
	   o_Energy_Bin_181      =>   energy_bin_neg_data(180 ),
	   o_Energy_Bin_182      =>   energy_bin_neg_data(181 ),
	   o_Energy_Bin_183      =>   energy_bin_neg_data(182 ),
	   o_Energy_Bin_184      =>   energy_bin_neg_data(183 ),
	   o_Energy_Bin_185      =>   energy_bin_neg_data(184 ),
	   o_Energy_Bin_186      =>   energy_bin_neg_data(185 ),
	   o_Energy_Bin_187      =>   energy_bin_neg_data(186 ),
	   o_Energy_Bin_188      =>   energy_bin_neg_data(187 ),
	   o_Energy_Bin_189      =>   energy_bin_neg_data(188 ),
	   o_Energy_Bin_190      =>   energy_bin_neg_data(189 ),
	   o_Energy_Bin_191      =>   energy_bin_neg_data(190 ),
	   o_Energy_Bin_192      =>   energy_bin_neg_data(191 ),
	   o_Energy_Bin_193      =>   energy_bin_neg_data(192 ),
	   o_Energy_Bin_194      =>   energy_bin_neg_data(193 ),
	   o_Energy_Bin_195      =>   energy_bin_neg_data(194 ),
	   o_Energy_Bin_196      =>   energy_bin_neg_data(195 ),
	   o_Energy_Bin_197      =>   energy_bin_neg_data(196 ),
	   o_Energy_Bin_198      =>   energy_bin_neg_data(197 ),
	   o_Energy_Bin_199      =>   energy_bin_neg_data(198 ),
	   o_Energy_Bin_200      =>   energy_bin_neg_data(199 ),
	   o_Energy_Bin_201      =>   energy_bin_neg_data(200 ),
	   o_Energy_Bin_202      =>   energy_bin_neg_data(201 ),
	   o_Energy_Bin_203      =>   energy_bin_neg_data(202 ),
	   o_Energy_Bin_204      =>   energy_bin_neg_data(203 ),
	   o_Energy_Bin_205      =>   energy_bin_neg_data(204 ),
	   o_Energy_Bin_206      =>   energy_bin_neg_data(205 ),
	   o_Energy_Bin_207      =>   energy_bin_neg_data(206 ),
	   o_Energy_Bin_208      =>   energy_bin_neg_data(207 ),
	   o_Energy_Bin_209      =>   energy_bin_neg_data(208 ),
	   o_Energy_Bin_210      =>   energy_bin_neg_data(209 ),
	   o_Energy_Bin_211      =>   energy_bin_neg_data(210 ),
	   o_Energy_Bin_212      =>   energy_bin_neg_data(211 ),
	   o_Energy_Bin_213      =>   energy_bin_neg_data(212 ),
	   o_Energy_Bin_214      =>   energy_bin_neg_data(213 ),
	   o_Energy_Bin_215      =>   energy_bin_neg_data(214 ),
	   o_Energy_Bin_216      =>   energy_bin_neg_data(215 ),
	   o_Energy_Bin_217      =>   energy_bin_neg_data(216 ),
	   o_Energy_Bin_218      =>   energy_bin_neg_data(217 ),
	   o_Energy_Bin_219      =>   energy_bin_neg_data(218 ),
	   o_Energy_Bin_220      =>   energy_bin_neg_data(219 ),
	   o_Energy_Bin_221      =>   energy_bin_neg_data(220 ),
	   o_Energy_Bin_222      =>   energy_bin_neg_data(221 ),
	   o_Energy_Bin_223      =>   energy_bin_neg_data(222 ),
	   o_Energy_Bin_224      =>   energy_bin_neg_data(223 ),
	   o_Energy_Bin_225      =>   energy_bin_neg_data(224 ),
	   o_Energy_Bin_226      =>   energy_bin_neg_data(225 ),
	   o_Energy_Bin_227      =>   energy_bin_neg_data(226 ),
	   o_Energy_Bin_228      =>   energy_bin_neg_data(227 ),
	   o_Energy_Bin_229      =>   energy_bin_neg_data(228 ),
	   o_Energy_Bin_230      =>   energy_bin_neg_data(229 ),
	   o_Energy_Bin_231      =>   energy_bin_neg_data(230 ),
	   o_Energy_Bin_232      =>   energy_bin_neg_data(231 ),
	   o_Energy_Bin_233      =>   energy_bin_neg_data(232 ),
	   o_Energy_Bin_234      =>   energy_bin_neg_data(233 ),
	   o_Energy_Bin_235      =>   energy_bin_neg_data(234 ),
	   o_Energy_Bin_236      =>   energy_bin_neg_data(235 ),
	   o_Energy_Bin_237      =>   energy_bin_neg_data(236 ),
	   o_Energy_Bin_238      =>   energy_bin_neg_data(237 ),
	   o_Energy_Bin_239      =>   energy_bin_neg_data(238 ),
	   o_Energy_Bin_240      =>   energy_bin_neg_data(239 ),
	   o_Energy_Bin_241      =>   energy_bin_neg_data(240 ),
	   o_Energy_Bin_242      =>   energy_bin_neg_data(241 ),
	   o_Energy_Bin_243      =>   energy_bin_neg_data(242 ),
	   o_Energy_Bin_244      =>   energy_bin_neg_data(243 ),
	   o_Energy_Bin_245      =>   energy_bin_neg_data(244 ),
	   o_Energy_Bin_246      =>   energy_bin_neg_data(245 ),
	   o_Energy_Bin_247      =>   energy_bin_neg_data(246 ),
	   o_Energy_Bin_248      =>   energy_bin_neg_data(247 ),
	   o_Energy_Bin_249      =>   energy_bin_neg_data(248 ),
	   o_Energy_Bin_250      =>   energy_bin_neg_data(249 ),
	   o_Energy_Bin_251      =>   energy_bin_neg_data(250 ),
	   o_Energy_Bin_252      =>   energy_bin_neg_data(251 ),
	   o_Energy_Bin_253      =>   energy_bin_neg_data(252 ),
	   o_Energy_Bin_254      =>   energy_bin_neg_data(253 ),
	   o_Energy_Bin_255      =>   energy_bin_neg_data(254 ),
	   o_Energy_Bin_256      =>   energy_bin_neg_data(255 ),
	   o_Energy_Bin_257      =>   energy_bin_neg_data(256 ),
	   o_Energy_Bin_258      =>   energy_bin_neg_data(257 ),
	   o_Energy_Bin_259      =>   energy_bin_neg_data(258 ),
	   o_Energy_Bin_260      =>   energy_bin_neg_data(259 ),
	   o_Energy_Bin_261      =>   energy_bin_neg_data(260 ),
	   o_Energy_Bin_262      =>   energy_bin_neg_data(261 ),
	   o_Energy_Bin_263      =>   energy_bin_neg_data(262 ),
	   o_Energy_Bin_264      =>   energy_bin_neg_data(263 ),
	   o_Energy_Bin_265      =>   energy_bin_neg_data(264 ),
	   o_Energy_Bin_266      =>   energy_bin_neg_data(265 ),
	   o_Energy_Bin_267      =>   energy_bin_neg_data(266 ),
	   o_Energy_Bin_268      =>   energy_bin_neg_data(267 ),
	   o_Energy_Bin_269      =>   energy_bin_neg_data(268 ),
	   o_Energy_Bin_270      =>   energy_bin_neg_data(269 ),
	   o_Energy_Bin_271      =>   energy_bin_neg_data(270 ),
	   o_Energy_Bin_272      =>   energy_bin_neg_data(271 ),
	   o_Energy_Bin_273      =>   energy_bin_neg_data(272 ),
	   o_Energy_Bin_274      =>   energy_bin_neg_data(273 ),
	   o_Energy_Bin_275      =>   energy_bin_neg_data(274 ),
	   o_Energy_Bin_276      =>   energy_bin_neg_data(275 ),
	   o_Energy_Bin_277      =>   energy_bin_neg_data(276 ),
	   o_Energy_Bin_278      =>   energy_bin_neg_data(277 ),
	   o_Energy_Bin_279      =>   energy_bin_neg_data(278 ),
	   o_Energy_Bin_280      =>   energy_bin_neg_data(279 ),
	   o_Energy_Bin_281      =>   energy_bin_neg_data(280 ),
	   o_Energy_Bin_282      =>   energy_bin_neg_data(281 ),
	   o_Energy_Bin_283      =>   energy_bin_neg_data(282 ),
	   o_Energy_Bin_284      =>   energy_bin_neg_data(283 ),
	   o_Energy_Bin_285      =>   energy_bin_neg_data(284 ),
	   o_Energy_Bin_286      =>   energy_bin_neg_data(285 ),
	   o_Energy_Bin_287      =>   energy_bin_neg_data(286 ),
	   o_Energy_Bin_288      =>   energy_bin_neg_data(287 ),
	   o_Energy_Bin_289      =>   energy_bin_neg_data(288 ),
	   o_Energy_Bin_290      =>   energy_bin_neg_data(289 ),
	   o_Energy_Bin_291      =>   energy_bin_neg_data(290 ),
	   o_Energy_Bin_292      =>   energy_bin_neg_data(291 ),
	   o_Energy_Bin_293      =>   energy_bin_neg_data(292 ),
	   o_Energy_Bin_294      =>   energy_bin_neg_data(293 ),
	   o_Energy_Bin_295      =>   energy_bin_neg_data(294 ),
	   o_Energy_Bin_296      =>   energy_bin_neg_data(295 ),
	   o_Energy_Bin_297      =>   energy_bin_neg_data(296 ),
	   o_Energy_Bin_298      =>   energy_bin_neg_data(297 ),
	   o_Energy_Bin_299      =>   energy_bin_neg_data(298 ),
	   o_Energy_Bin_300      =>   energy_bin_neg_data(299 ),
	   o_Energy_Bin_301      =>   energy_bin_neg_data(300 ),
	   o_Energy_Bin_302      =>   energy_bin_neg_data(301 ),
	   o_Energy_Bin_303      =>   energy_bin_neg_data(302 ),
	   o_Energy_Bin_304      =>   energy_bin_neg_data(303 ),
	   o_Energy_Bin_305      =>   energy_bin_neg_data(304 ),
	   o_Energy_Bin_306      =>   energy_bin_neg_data(305 ),
	   o_Energy_Bin_307      =>   energy_bin_neg_data(306 ),
	   o_Energy_Bin_308      =>   energy_bin_neg_data(307 ),
	   o_Energy_Bin_309      =>   energy_bin_neg_data(308 ),
	   o_Energy_Bin_310      =>   energy_bin_neg_data(309 ),
	   o_Energy_Bin_311      =>   energy_bin_neg_data(310 ),
	   o_Energy_Bin_312      =>   energy_bin_neg_data(311 ),
	   o_Energy_Bin_313      =>   energy_bin_neg_data(312 ),
	   o_Energy_Bin_314      =>   energy_bin_neg_data(313 ),
	   o_Energy_Bin_315      =>   energy_bin_neg_data(314 ),
	   o_Energy_Bin_316      =>   energy_bin_neg_data(315 ),
	   o_Energy_Bin_317      =>   energy_bin_neg_data(316 ),
	   o_Energy_Bin_318      =>   energy_bin_neg_data(317 ),
	   o_Energy_Bin_319      =>   energy_bin_neg_data(318 ),
	   o_Energy_Bin_320      =>   energy_bin_neg_data(319 ),
	   o_Energy_Bin_321      =>   energy_bin_neg_data(320 ),
	   o_Energy_Bin_322      =>   energy_bin_neg_data(321 ),
	   o_Energy_Bin_323      =>   energy_bin_neg_data(322 ),
	   o_Energy_Bin_324      =>   energy_bin_neg_data(323 ),
	   o_Energy_Bin_325      =>   energy_bin_neg_data(324 ),
	   o_Energy_Bin_326      =>   energy_bin_neg_data(325 ),
	   o_Energy_Bin_327      =>   energy_bin_neg_data(326 ),
	   o_Energy_Bin_328      =>   energy_bin_neg_data(327 ),
	   o_Energy_Bin_329      =>   energy_bin_neg_data(328 ),
	   o_Energy_Bin_330      =>   energy_bin_neg_data(329 ),
	   o_Energy_Bin_331      =>   energy_bin_neg_data(330 ),
	   o_Energy_Bin_332      =>   energy_bin_neg_data(331 ),
	   o_Energy_Bin_333      =>   energy_bin_neg_data(332 ),
	   o_Energy_Bin_334      =>   energy_bin_neg_data(333 ),
	   o_Energy_Bin_335      =>   energy_bin_neg_data(334 ),
	   o_Energy_Bin_336      =>   energy_bin_neg_data(335 ),
	   o_Energy_Bin_337      =>   energy_bin_neg_data(336 ),
	   o_Energy_Bin_338      =>   energy_bin_neg_data(337 ),
	   o_Energy_Bin_339      =>   energy_bin_neg_data(338 ),
	   o_Energy_Bin_340      =>   energy_bin_neg_data(339 ),
	   o_Energy_Bin_341      =>   energy_bin_neg_data(340 ),
	   o_Energy_Bin_342      =>   energy_bin_neg_data(341 ),
	   o_Energy_Bin_343      =>   energy_bin_neg_data(342 ),
	   o_Energy_Bin_344      =>   energy_bin_neg_data(343 ),
	   o_Energy_Bin_345      =>   energy_bin_neg_data(344 ),
	   o_Energy_Bin_346      =>   energy_bin_neg_data(345 ),
	   o_Energy_Bin_347      =>   energy_bin_neg_data(346 ),
	   o_Energy_Bin_348      =>   energy_bin_neg_data(347 ),
	   o_Energy_Bin_349      =>   energy_bin_neg_data(348 ),
	   o_Energy_Bin_350      =>   energy_bin_neg_data(349 ),
	   o_Energy_Bin_351      =>   energy_bin_neg_data(350 ),
	   o_Energy_Bin_352      =>   energy_bin_neg_data(351 ),
	   o_Energy_Bin_353      =>   energy_bin_neg_data(352 ),
	   o_Energy_Bin_354      =>   energy_bin_neg_data(353 ),
	   o_Energy_Bin_355      =>   energy_bin_neg_data(354 ),
	   o_Energy_Bin_356      =>   energy_bin_neg_data(355 ),
	   o_Energy_Bin_357      =>   energy_bin_neg_data(356 ),
	   o_Energy_Bin_358      =>   energy_bin_neg_data(357 ),
	   o_Energy_Bin_359      =>   energy_bin_neg_data(358 ),
	   o_Energy_Bin_360      =>   energy_bin_neg_data(359 ),
	   o_Energy_Bin_361      =>   energy_bin_neg_data(360 ),
	   o_Energy_Bin_362      =>   energy_bin_neg_data(361 ),
	   o_Energy_Bin_363      =>   energy_bin_neg_data(362 ),
	   o_Energy_Bin_364      =>   energy_bin_neg_data(363 ),
	   o_Energy_Bin_365      =>   energy_bin_neg_data(364 ),
	   o_Energy_Bin_366      =>   energy_bin_neg_data(365 ),
	   o_Energy_Bin_367      =>   energy_bin_neg_data(366 ),
	   o_Energy_Bin_368      =>   energy_bin_neg_data(367 ),
	   o_Energy_Bin_369      =>   energy_bin_neg_data(368 ),
	   o_Energy_Bin_370      =>   energy_bin_neg_data(369 ),
	   o_Energy_Bin_371      =>   energy_bin_neg_data(370 ),
	   o_Energy_Bin_372      =>   energy_bin_neg_data(371 ),
	   o_Energy_Bin_373      =>   energy_bin_neg_data(372 ),
	   o_Energy_Bin_374      =>   energy_bin_neg_data(373 ),
	   o_Energy_Bin_375      =>   energy_bin_neg_data(374 ),
	   o_Energy_Bin_376      =>   energy_bin_neg_data(375 ),
	   o_Energy_Bin_377      =>   energy_bin_neg_data(376 ),
	   o_Energy_Bin_378      =>   energy_bin_neg_data(377 ),
	   o_Energy_Bin_379      =>   energy_bin_neg_data(378 ),
	   o_Energy_Bin_380      =>   energy_bin_neg_data(379 ),
	   o_Energy_Bin_381      =>   energy_bin_neg_data(380 ),
	   o_Energy_Bin_382      =>   energy_bin_neg_data(381 ),
	   o_Energy_Bin_383      =>   energy_bin_neg_data(382 ),
	   o_Energy_Bin_384      =>   energy_bin_neg_data(383 ),
	   o_Energy_Bin_385      =>   energy_bin_neg_data(384 ),
	   o_Energy_Bin_386      =>   energy_bin_neg_data(385 ),
	   o_Energy_Bin_387      =>   energy_bin_neg_data(386 ),
	   o_Energy_Bin_388      =>   energy_bin_neg_data(387 ),
	   o_Energy_Bin_389      =>   energy_bin_neg_data(388 ),
	   o_Energy_Bin_390      =>   energy_bin_neg_data(389 ),
	   o_Energy_Bin_391      =>   energy_bin_neg_data(390 ),
	   o_Energy_Bin_392      =>   energy_bin_neg_data(391 ),
	   o_Energy_Bin_393      =>   energy_bin_neg_data(392 ),
	   o_Energy_Bin_394      =>   energy_bin_neg_data(393 ),
	   o_Energy_Bin_395      =>   energy_bin_neg_data(394 ),
	   o_Energy_Bin_396      =>   energy_bin_neg_data(395 ),
	   o_Energy_Bin_397      =>   energy_bin_neg_data(396 ),
	   o_Energy_Bin_398      =>   energy_bin_neg_data(397 ),
	   o_Energy_Bin_399      =>   energy_bin_neg_data(398 ),
	   o_Energy_Bin_400      =>   energy_bin_neg_data(399 ),
	   o_Energy_Bin_401      =>   energy_bin_neg_data(400 ),
	   o_Energy_Bin_402      =>   energy_bin_neg_data(401 ),
	   o_Energy_Bin_403      =>   energy_bin_neg_data(402 ),
	   o_Energy_Bin_404      =>   energy_bin_neg_data(403 ),
	   o_Energy_Bin_405      =>   energy_bin_neg_data(404 ),
	   o_Energy_Bin_406      =>   energy_bin_neg_data(405 ),
	   o_Energy_Bin_407      =>   energy_bin_neg_data(406 ),
	   o_Energy_Bin_408      =>   energy_bin_neg_data(407 ),
	   o_Energy_Bin_409      =>   energy_bin_neg_data(408 ),
	   o_Energy_Bin_410      =>   energy_bin_neg_data(409 ),
	   o_Energy_Bin_411      =>   energy_bin_neg_data(410 ),
	   o_Energy_Bin_412      =>   energy_bin_neg_data(411 ),
	   o_Energy_Bin_413      =>   energy_bin_neg_data(412 ),
	   o_Energy_Bin_414      =>   energy_bin_neg_data(413 ),
	   o_Energy_Bin_415      =>   energy_bin_neg_data(414 ),
	   o_Energy_Bin_416      =>   energy_bin_neg_data(415 ),
	   o_Energy_Bin_417      =>   energy_bin_neg_data(416 ),
	   o_Energy_Bin_418      =>   energy_bin_neg_data(417 ),
	   o_Energy_Bin_419      =>   energy_bin_neg_data(418 ),
	   o_Energy_Bin_420      =>   energy_bin_neg_data(419 ),
	   o_Energy_Bin_421      =>   energy_bin_neg_data(420 ),
	   o_Energy_Bin_422      =>   energy_bin_neg_data(421 ),
	   o_Energy_Bin_423      =>   energy_bin_neg_data(422 ),
	   o_Energy_Bin_424      =>   energy_bin_neg_data(423 ),
	   o_Energy_Bin_425      =>   energy_bin_neg_data(424 ),
	   o_Energy_Bin_426      =>   energy_bin_neg_data(425 ),
	   o_Energy_Bin_427      =>   energy_bin_neg_data(426 ),
	   o_Energy_Bin_428      =>   energy_bin_neg_data(427 ),
	   o_Energy_Bin_429      =>   energy_bin_neg_data(428 ),
	   o_Energy_Bin_430      =>   energy_bin_neg_data(429 ),
	   o_Energy_Bin_431      =>   energy_bin_neg_data(430 ),
	   o_Energy_Bin_432      =>   energy_bin_neg_data(431 ),
	   o_Energy_Bin_433      =>   energy_bin_neg_data(432 ),
	   o_Energy_Bin_434      =>   energy_bin_neg_data(433 ),
	   o_Energy_Bin_435      =>   energy_bin_neg_data(434 ),
	   o_Energy_Bin_436      =>   energy_bin_neg_data(435 ),
	   o_Energy_Bin_437      =>   energy_bin_neg_data(436 ),
	   o_Energy_Bin_438      =>   energy_bin_neg_data(437 ),
	   o_Energy_Bin_439      =>   energy_bin_neg_data(438 ),
	   o_Energy_Bin_440      =>   energy_bin_neg_data(439 ),
	   o_Energy_Bin_441      =>   energy_bin_neg_data(440 ),
	   o_Energy_Bin_442      =>   energy_bin_neg_data(441 ),
	   o_Energy_Bin_443      =>   energy_bin_neg_data(442 ),
	   o_Energy_Bin_444      =>   energy_bin_neg_data(443 ),
	   o_Energy_Bin_445      =>   energy_bin_neg_data(444 ),
	   o_Energy_Bin_446      =>   energy_bin_neg_data(445 ),
	   o_Energy_Bin_447      =>   energy_bin_neg_data(446 ),
	   o_Energy_Bin_448      =>   energy_bin_neg_data(447 ),
	   o_Energy_Bin_449      =>   energy_bin_neg_data(448 ),
	   o_Energy_Bin_450      =>   energy_bin_neg_data(449 ),
	   o_Energy_Bin_451      =>   energy_bin_neg_data(450 ),
	   o_Energy_Bin_452      =>   energy_bin_neg_data(451 ),
	   o_Energy_Bin_453      =>   energy_bin_neg_data(452 ),
	   o_Energy_Bin_454      =>   energy_bin_neg_data(453 ),
	   o_Energy_Bin_455      =>   energy_bin_neg_data(454 ),
	   o_Energy_Bin_456      =>   energy_bin_neg_data(455 ),
	   o_Energy_Bin_457      =>   energy_bin_neg_data(456 ),
	   o_Energy_Bin_458      =>   energy_bin_neg_data(457 ),
	   o_Energy_Bin_459      =>   energy_bin_neg_data(458 ),
	   o_Energy_Bin_460      =>   energy_bin_neg_data(459 ),
	   o_Energy_Bin_461      =>   energy_bin_neg_data(460 ),
	   o_Energy_Bin_462      =>   energy_bin_neg_data(461 ),
	   o_Energy_Bin_463      =>   energy_bin_neg_data(462 ),
	   o_Energy_Bin_464      =>   energy_bin_neg_data(463 ),
	   o_Energy_Bin_465      =>   energy_bin_neg_data(464 ),
	   o_Energy_Bin_466      =>   energy_bin_neg_data(465 ),
	   o_Energy_Bin_467      =>   energy_bin_neg_data(466 ),
	   o_Energy_Bin_468      =>   energy_bin_neg_data(467 ),
	   o_Energy_Bin_469      =>   energy_bin_neg_data(468 ),
	   o_Energy_Bin_470      =>   energy_bin_neg_data(469 ),
	   o_Energy_Bin_471      =>   energy_bin_neg_data(470 ),
	   o_Energy_Bin_472      =>   energy_bin_neg_data(471 ),
	   o_Energy_Bin_473      =>   energy_bin_neg_data(472 ),
	   o_Energy_Bin_474      =>   energy_bin_neg_data(473 ),
	   o_Energy_Bin_475      =>   energy_bin_neg_data(474 ),
	   o_Energy_Bin_476      =>   energy_bin_neg_data(475 ),
	   o_Energy_Bin_477      =>   energy_bin_neg_data(476 ),
	   o_Energy_Bin_478      =>   energy_bin_neg_data(477 ),
	   o_Energy_Bin_479      =>   energy_bin_neg_data(478 ),
	   o_Energy_Bin_480      =>   energy_bin_neg_data(479 ),
	   o_Energy_Bin_481      =>   energy_bin_neg_data(480 ),
	   o_Energy_Bin_482      =>   energy_bin_neg_data(481 ),
	   o_Energy_Bin_483      =>   energy_bin_neg_data(482 ),
	   o_Energy_Bin_484      =>   energy_bin_neg_data(483 ),
	   o_Energy_Bin_485      =>   energy_bin_neg_data(484 ),
	   o_Energy_Bin_486      =>   energy_bin_neg_data(485 ),
	   o_Energy_Bin_487      =>   energy_bin_neg_data(486 ),
	   o_Energy_Bin_488      =>   energy_bin_neg_data(487 ),
	   o_Energy_Bin_489      =>   energy_bin_neg_data(488 ),
	   o_Energy_Bin_490      =>   energy_bin_neg_data(489 ),
	   o_Energy_Bin_491      =>   energy_bin_neg_data(490 ),
	   o_Energy_Bin_492      =>   energy_bin_neg_data(491 ),
	   o_Energy_Bin_493      =>   energy_bin_neg_data(492 ),
	   o_Energy_Bin_494      =>   energy_bin_neg_data(493 ),
	   o_Energy_Bin_495      =>   energy_bin_neg_data(494 ),
	   o_Energy_Bin_496      =>   energy_bin_neg_data(495 ),
	   o_Energy_Bin_497      =>   energy_bin_neg_data(496 ),
	   o_Energy_Bin_498      =>   energy_bin_neg_data(497 ),
	   o_Energy_Bin_499      =>   energy_bin_neg_data(498 ),
	   o_Energy_Bin_500      =>   energy_bin_neg_data(499 ),
	   o_Energy_Bin_501      =>   energy_bin_neg_data(500 ),
	   o_Energy_Bin_502      =>   energy_bin_neg_data(501 ),
	   o_Energy_Bin_503      =>   energy_bin_neg_data(502 ),
	   o_Energy_Bin_504      =>   energy_bin_neg_data(503 ),
	   o_Energy_Bin_505      =>   energy_bin_neg_data(504 ),
	   o_Energy_Bin_506      =>   energy_bin_neg_data(505 ),
	   o_Energy_Bin_507      =>   energy_bin_neg_data(506 ),
	   o_Energy_Bin_508      =>   energy_bin_neg_data(507 ),
	   o_Energy_Bin_509      =>   energy_bin_neg_data(508 ),
	   o_Energy_Bin_510      =>   energy_bin_neg_data(509 ),
	   o_Energy_Bin_511      =>   energy_bin_neg_data(510 ),
	   o_Energy_Bin_512      =>   energy_bin_neg_data(511 ),
	   o_Energy_Bin_513      =>   energy_bin_neg_data(512 ),
	   o_Energy_Bin_514      =>   energy_bin_neg_data(513 ),
	   o_Energy_Bin_515      =>   energy_bin_neg_data(514 ),
	   o_Energy_Bin_516      =>   energy_bin_neg_data(515 ),
	   o_Energy_Bin_517      =>   energy_bin_neg_data(516 ),
	   o_Energy_Bin_518      =>   energy_bin_neg_data(517 ),
	   o_Energy_Bin_519      =>   energy_bin_neg_data(518 ),
	   o_Energy_Bin_520      =>   energy_bin_neg_data(519 ),
	   o_Energy_Bin_521      =>   energy_bin_neg_data(520 ),
	   o_Energy_Bin_522      =>   energy_bin_neg_data(521 ),
	   o_Energy_Bin_523      =>   energy_bin_neg_data(522 ),
	   o_Energy_Bin_524      =>   energy_bin_neg_data(523 ),
	   o_Energy_Bin_525      =>   energy_bin_neg_data(524 ),
	   o_Energy_Bin_526      =>   energy_bin_neg_data(525 ),
	   o_Energy_Bin_527      =>   energy_bin_neg_data(526 ),
	   o_Energy_Bin_528      =>   energy_bin_neg_data(527 ),
	   o_Energy_Bin_529      =>   energy_bin_neg_data(528 ),
	   o_Energy_Bin_530      =>   energy_bin_neg_data(529 ),
	   o_Energy_Bin_531      =>   energy_bin_neg_data(530 ),
	   o_Energy_Bin_532      =>   energy_bin_neg_data(531 ),
	   o_Energy_Bin_533      =>   energy_bin_neg_data(532 ),
	   o_Energy_Bin_534      =>   energy_bin_neg_data(533 ),
	   o_Energy_Bin_535      =>   energy_bin_neg_data(534 ),
	   o_Energy_Bin_536      =>   energy_bin_neg_data(535 ),
	   o_Energy_Bin_537      =>   energy_bin_neg_data(536 ),
	   o_Energy_Bin_538      =>   energy_bin_neg_data(537 ),
	   o_Energy_Bin_539      =>   energy_bin_neg_data(538 ),
	   o_Energy_Bin_540      =>   energy_bin_neg_data(539 ),
	   o_Energy_Bin_541      =>   energy_bin_neg_data(540 ),
	   o_Energy_Bin_542      =>   energy_bin_neg_data(541 ),
	   o_Energy_Bin_543      =>   energy_bin_neg_data(542 ),
	   o_Energy_Bin_544      =>   energy_bin_neg_data(543 ),
	   o_Energy_Bin_545      =>   energy_bin_neg_data(544 ),
	   o_Energy_Bin_546      =>   energy_bin_neg_data(545 ),
	   o_Energy_Bin_547      =>   energy_bin_neg_data(546 ),
	   o_Energy_Bin_548      =>   energy_bin_neg_data(547 ),
	   o_Energy_Bin_549      =>   energy_bin_neg_data(548 ),
	   o_Energy_Bin_550      =>   energy_bin_neg_data(549 ),
	   o_Energy_Bin_551      =>   energy_bin_neg_data(550 ),
	   o_Energy_Bin_552      =>   energy_bin_neg_data(551 ),
	   o_Energy_Bin_553      =>   energy_bin_neg_data(552 ),
	   o_Energy_Bin_554      =>   energy_bin_neg_data(553 ),
	   o_Energy_Bin_555      =>   energy_bin_neg_data(554 ),
	   o_Energy_Bin_556      =>   energy_bin_neg_data(555 ),
	   o_Energy_Bin_557      =>   energy_bin_neg_data(556 ),
	   o_Energy_Bin_558      =>   energy_bin_neg_data(557 ),
	   o_Energy_Bin_559      =>   energy_bin_neg_data(558 ),
	   o_Energy_Bin_560      =>   energy_bin_neg_data(559 ),
	   o_Energy_Bin_561      =>   energy_bin_neg_data(560 ),
	   o_Energy_Bin_562      =>   energy_bin_neg_data(561 ),
	   o_Energy_Bin_563      =>   energy_bin_neg_data(562 ),
	   o_Energy_Bin_564      =>   energy_bin_neg_data(563 ),
	   o_Energy_Bin_565      =>   energy_bin_neg_data(564 ),
	   o_Energy_Bin_566      =>   energy_bin_neg_data(565 ),
	   o_Energy_Bin_567      =>   energy_bin_neg_data(566 ),
	   o_Energy_Bin_568      =>   energy_bin_neg_data(567 ),
	   o_Energy_Bin_569      =>   energy_bin_neg_data(568 ),
	   o_Energy_Bin_570      =>   energy_bin_neg_data(569 ),
	   o_Energy_Bin_571      =>   energy_bin_neg_data(570 ),
	   o_Energy_Bin_572      =>   energy_bin_neg_data(571 ),
	   o_Energy_Bin_573      =>   energy_bin_neg_data(572 ),
	   o_Energy_Bin_574      =>   energy_bin_neg_data(573 ),
	   o_Energy_Bin_575      =>   energy_bin_neg_data(574 ),
	   o_Energy_Bin_576      =>   energy_bin_neg_data(575 ),
	   o_Energy_Bin_577      =>   energy_bin_neg_data(576 ),
	   o_Energy_Bin_578      =>   energy_bin_neg_data(577 ),
	   o_Energy_Bin_579      =>   energy_bin_neg_data(578 ),
	   o_Energy_Bin_580      =>   energy_bin_neg_data(579 ),
	   o_Energy_Bin_581      =>   energy_bin_neg_data(580 ),
	   o_Energy_Bin_582      =>   energy_bin_neg_data(581 ),
	   o_Energy_Bin_583      =>   energy_bin_neg_data(582 ),
	   o_Energy_Bin_584      =>   energy_bin_neg_data(583 ),
	   o_Energy_Bin_585      =>   energy_bin_neg_data(584 ),
	   o_Energy_Bin_586      =>   energy_bin_neg_data(585 ),
	   o_Energy_Bin_587      =>   energy_bin_neg_data(586 ),
	   o_Energy_Bin_588      =>   energy_bin_neg_data(587 ),
	   o_Energy_Bin_589      =>   energy_bin_neg_data(588 ),
	   o_Energy_Bin_590      =>   energy_bin_neg_data(589 ),
	   o_Energy_Bin_591      =>   energy_bin_neg_data(590 ),
	   o_Energy_Bin_592      =>   energy_bin_neg_data(591 ),
	   o_Energy_Bin_593      =>   energy_bin_neg_data(592 ),
	   o_Energy_Bin_594      =>   energy_bin_neg_data(593 ),
	   o_Energy_Bin_595      =>   energy_bin_neg_data(594 ),
	   o_Energy_Bin_596      =>   energy_bin_neg_data(595 ),
	   o_Energy_Bin_597      =>   energy_bin_neg_data(596 ),
	   o_Energy_Bin_598      =>   energy_bin_neg_data(597 ),
	   o_Energy_Bin_599      =>   energy_bin_neg_data(598 ),
	   o_Energy_Bin_600      =>   energy_bin_neg_data(599 ),
	   o_Energy_Bin_601      =>   energy_bin_neg_data(600 ),
	   o_Energy_Bin_602      =>   energy_bin_neg_data(601 ),
	   o_Energy_Bin_603      =>   energy_bin_neg_data(602 ),
	   o_Energy_Bin_604      =>   energy_bin_neg_data(603 ),
	   o_Energy_Bin_605      =>   energy_bin_neg_data(604 ),
	   o_Energy_Bin_606      =>   energy_bin_neg_data(605 ),
	   o_Energy_Bin_607      =>   energy_bin_neg_data(606 ),
	   o_Energy_Bin_608      =>   energy_bin_neg_data(607 ),
	   o_Energy_Bin_609      =>   energy_bin_neg_data(608 ),
	   o_Energy_Bin_610      =>   energy_bin_neg_data(609 ),
	   o_Energy_Bin_611      =>   energy_bin_neg_data(610 ),
	   o_Energy_Bin_612      =>   energy_bin_neg_data(611 ),
	   o_Energy_Bin_613      =>   energy_bin_neg_data(612 ),
	   o_Energy_Bin_614      =>   energy_bin_neg_data(613 ),
	   o_Energy_Bin_615      =>   energy_bin_neg_data(614 ),
	   o_Energy_Bin_616      =>   energy_bin_neg_data(615 ),
	   o_Energy_Bin_617      =>   energy_bin_neg_data(616 ),
	   o_Energy_Bin_618      =>   energy_bin_neg_data(617 ),
	   o_Energy_Bin_619      =>   energy_bin_neg_data(618 ),
	   o_Energy_Bin_620      =>   energy_bin_neg_data(619 ),
	   o_Energy_Bin_621      =>   energy_bin_neg_data(620 ),
	   o_Energy_Bin_622      =>   energy_bin_neg_data(621 ),
	   o_Energy_Bin_623      =>   energy_bin_neg_data(622 ),
	   o_Energy_Bin_624      =>   energy_bin_neg_data(623 ),
	   o_Energy_Bin_625      =>   energy_bin_neg_data(624 ),
	   o_Energy_Bin_626      =>   energy_bin_neg_data(625 ),
	   o_Energy_Bin_627      =>   energy_bin_neg_data(626 ),
	   o_Energy_Bin_628      =>   energy_bin_neg_data(627 ),
	   o_Energy_Bin_629      =>   energy_bin_neg_data(628 ),
	   o_Energy_Bin_630      =>   energy_bin_neg_data(629 ),
	   o_Energy_Bin_631      =>   energy_bin_neg_data(630 ),
	   o_Energy_Bin_632      =>   energy_bin_neg_data(631 ),
	   o_Energy_Bin_633      =>   energy_bin_neg_data(632 ),
	   o_Energy_Bin_634      =>   energy_bin_neg_data(633 ),
	   o_Energy_Bin_635      =>   energy_bin_neg_data(634 ),
	   o_Energy_Bin_636      =>   energy_bin_neg_data(635 ),
	   o_Energy_Bin_637      =>   energy_bin_neg_data(636 ),
	   o_Energy_Bin_638      =>   energy_bin_neg_data(637 ),
	   o_Energy_Bin_639      =>   energy_bin_neg_data(638 ),
	   o_Energy_Bin_640      =>   energy_bin_neg_data(639 ),
	   o_Energy_Bin_641      =>   energy_bin_neg_data(640 ),
	   o_Energy_Bin_642      =>   energy_bin_neg_data(641 ),
	   o_Energy_Bin_643      =>   energy_bin_neg_data(642 ),
	   o_Energy_Bin_644      =>   energy_bin_neg_data(643 ),
	   o_Energy_Bin_645      =>   energy_bin_neg_data(644 ),
	   o_Energy_Bin_646      =>   energy_bin_neg_data(645 ),
	   o_Energy_Bin_647      =>   energy_bin_neg_data(646 ),
	   o_Energy_Bin_648      =>   energy_bin_neg_data(647 ),
	   o_Energy_Bin_649      =>   energy_bin_neg_data(648 ),
	   o_Energy_Bin_650      =>   energy_bin_neg_data(649 ),
	   o_Energy_Bin_651      =>   energy_bin_neg_data(650 ),
	   o_Energy_Bin_652      =>   energy_bin_neg_data(651 ),
	   o_Energy_Bin_653      =>   energy_bin_neg_data(652 ),
	   o_Energy_Bin_654      =>   energy_bin_neg_data(653 ),
	   o_Energy_Bin_655      =>   energy_bin_neg_data(654 ),
	   o_Energy_Bin_656      =>   energy_bin_neg_data(655 ),
	   o_Energy_Bin_657      =>   energy_bin_neg_data(656 ),
	   o_Energy_Bin_658      =>   energy_bin_neg_data(657 ),
	   o_Energy_Bin_659      =>   energy_bin_neg_data(658 ),
	   o_Energy_Bin_660      =>   energy_bin_neg_data(659 ),
	   o_Energy_Bin_661      =>   energy_bin_neg_data(660 ),
	   o_Energy_Bin_662      =>   energy_bin_neg_data(661 ),
	   o_Energy_Bin_663      =>   energy_bin_neg_data(662 ),
	   o_Energy_Bin_664      =>   energy_bin_neg_data(663 ),
	   o_Energy_Bin_665      =>   energy_bin_neg_data(664 ),
	   o_Energy_Bin_666      =>   energy_bin_neg_data(665 ),
	   o_Energy_Bin_667      =>   energy_bin_neg_data(666 ),
	   o_Energy_Bin_668      =>   energy_bin_neg_data(667 ),
	   o_Energy_Bin_669      =>   energy_bin_neg_data(668 ),
	   o_Energy_Bin_670      =>   energy_bin_neg_data(669 ),
	   o_Energy_Bin_671      =>   energy_bin_neg_data(670 ),
	   o_Energy_Bin_672      =>   energy_bin_neg_data(671 ),
	   o_Energy_Bin_673      =>   energy_bin_neg_data(672 ),
	   o_Energy_Bin_674      =>   energy_bin_neg_data(673 ),
	   o_Energy_Bin_675      =>   energy_bin_neg_data(674 ),
	   o_Energy_Bin_676      =>   energy_bin_neg_data(675 ),
	   o_Energy_Bin_677      =>   energy_bin_neg_data(676 ),
	   o_Energy_Bin_678      =>   energy_bin_neg_data(677 ),
	   o_Energy_Bin_679      =>   energy_bin_neg_data(678 ),
	   o_Energy_Bin_680      =>   energy_bin_neg_data(679 ),
	   o_Energy_Bin_681      =>   energy_bin_neg_data(680 ),
	   o_Energy_Bin_682      =>   energy_bin_neg_data(681 ),
	   o_Energy_Bin_683      =>   energy_bin_neg_data(682 ),
	   o_Energy_Bin_684      =>   energy_bin_neg_data(683 ),
	   o_Energy_Bin_685      =>   energy_bin_neg_data(684 ),
	   o_Energy_Bin_686      =>   energy_bin_neg_data(685 ),
	   o_Energy_Bin_687      =>   energy_bin_neg_data(686 ),
	   o_Energy_Bin_688      =>   energy_bin_neg_data(687 ),
	   o_Energy_Bin_689      =>   energy_bin_neg_data(688 ),
	   o_Energy_Bin_690      =>   energy_bin_neg_data(689 ),
	   o_Energy_Bin_691      =>   energy_bin_neg_data(690 ),
	   o_Energy_Bin_692      =>   energy_bin_neg_data(691 ),
	   o_Energy_Bin_693      =>   energy_bin_neg_data(692 ),
	   o_Energy_Bin_694      =>   energy_bin_neg_data(693 ),
	   o_Energy_Bin_695      =>   energy_bin_neg_data(694 ),
	   o_Energy_Bin_696      =>   energy_bin_neg_data(695 ),
	   o_Energy_Bin_697      =>   energy_bin_neg_data(696 ),
	   o_Energy_Bin_698      =>   energy_bin_neg_data(697 ),
	   o_Energy_Bin_699      =>   energy_bin_neg_data(698 ),
	   o_Energy_Bin_700      =>   energy_bin_neg_data(699 ),
	   o_Energy_Bin_701      =>   energy_bin_neg_data(700 ),
	   o_Energy_Bin_702      =>   energy_bin_neg_data(701 ),
	   o_Energy_Bin_703      =>   energy_bin_neg_data(702 ),
	   o_Energy_Bin_704      =>   energy_bin_neg_data(703 ),
	   o_Energy_Bin_705      =>   energy_bin_neg_data(704 ),
	   o_Energy_Bin_706      =>   energy_bin_neg_data(705 ),
	   o_Energy_Bin_707      =>   energy_bin_neg_data(706 ),
	   o_Energy_Bin_708      =>   energy_bin_neg_data(707 ),
	   o_Energy_Bin_709      =>   energy_bin_neg_data(708 ),
	   o_Energy_Bin_710      =>   energy_bin_neg_data(709 ),
	   o_Energy_Bin_711      =>   energy_bin_neg_data(710 ),
	   o_Energy_Bin_712      =>   energy_bin_neg_data(711 ),
	   o_Energy_Bin_713      =>   energy_bin_neg_data(712 ),
	   o_Energy_Bin_714      =>   energy_bin_neg_data(713 ),
	   o_Energy_Bin_715      =>   energy_bin_neg_data(714 ),
	   o_Energy_Bin_716      =>   energy_bin_neg_data(715 ),
	   o_Energy_Bin_717      =>   energy_bin_neg_data(716 ),
	   o_Energy_Bin_718      =>   energy_bin_neg_data(717 ),
	   o_Energy_Bin_719      =>   energy_bin_neg_data(718 ),
	   o_Energy_Bin_720      =>   energy_bin_neg_data(719 ),
	   o_Energy_Bin_721      =>   energy_bin_neg_data(720 ),
	   o_Energy_Bin_722      =>   energy_bin_neg_data(721 ),
	   o_Energy_Bin_723      =>   energy_bin_neg_data(722 ),
	   o_Energy_Bin_724      =>   energy_bin_neg_data(723 ),
	   o_Energy_Bin_725      =>   energy_bin_neg_data(724 ),
	   o_Energy_Bin_726      =>   energy_bin_neg_data(725 ),
	   o_Energy_Bin_727      =>   energy_bin_neg_data(726 ),
	   o_Energy_Bin_728      =>   energy_bin_neg_data(727 ),
	   o_Energy_Bin_729      =>   energy_bin_neg_data(728 ),
	   o_Energy_Bin_730      =>   energy_bin_neg_data(729 ),
	   o_Energy_Bin_731      =>   energy_bin_neg_data(730 ),
	   o_Energy_Bin_732      =>   energy_bin_neg_data(731 ),
	   o_Energy_Bin_733      =>   energy_bin_neg_data(732 ),
	   o_Energy_Bin_734      =>   energy_bin_neg_data(733 ),
	   o_Energy_Bin_735      =>   energy_bin_neg_data(734 ),
	   o_Energy_Bin_736      =>   energy_bin_neg_data(735 ),
	   o_Energy_Bin_737      =>   energy_bin_neg_data(736 ),
	   o_Energy_Bin_738      =>   energy_bin_neg_data(737 ),
	   o_Energy_Bin_739      =>   energy_bin_neg_data(738 ),
	   o_Energy_Bin_740      =>   energy_bin_neg_data(739 ),
	   o_Energy_Bin_741      =>   energy_bin_neg_data(740 ),
	   o_Energy_Bin_742      =>   energy_bin_neg_data(741 ),
	   o_Energy_Bin_743      =>   energy_bin_neg_data(742 ),
	   o_Energy_Bin_744      =>   energy_bin_neg_data(743 ),
	   o_Energy_Bin_745      =>   energy_bin_neg_data(744 ),
	   o_Energy_Bin_746      =>   energy_bin_neg_data(745 ),
	   o_Energy_Bin_747      =>   energy_bin_neg_data(746 ),
	   o_Energy_Bin_748      =>   energy_bin_neg_data(747 ),
	   o_Energy_Bin_749      =>   energy_bin_neg_data(748 ),
	   o_Energy_Bin_750      =>   energy_bin_neg_data(749 ),
	   o_Energy_Bin_751      =>   energy_bin_neg_data(750 ),
	   o_Energy_Bin_752      =>   energy_bin_neg_data(751 ),
	   o_Energy_Bin_753      =>   energy_bin_neg_data(752 ),
	   o_Energy_Bin_754      =>   energy_bin_neg_data(753 ),
	   o_Energy_Bin_755      =>   energy_bin_neg_data(754 ),
	   o_Energy_Bin_756      =>   energy_bin_neg_data(755 ),
	   o_Energy_Bin_757      =>   energy_bin_neg_data(756 ),
	   o_Energy_Bin_758      =>   energy_bin_neg_data(757 ),
	   o_Energy_Bin_759      =>   energy_bin_neg_data(758 ),
	   o_Energy_Bin_760      =>   energy_bin_neg_data(759 ),
	   o_Energy_Bin_761      =>   energy_bin_neg_data(760 ),
	   o_Energy_Bin_762      =>   energy_bin_neg_data(761 ),
	   o_Energy_Bin_763      =>   energy_bin_neg_data(762 ),
	   o_Energy_Bin_764      =>   energy_bin_neg_data(763 ),
	   o_Energy_Bin_765      =>   energy_bin_neg_data(764 ),
	   o_Energy_Bin_766      =>   energy_bin_neg_data(765 ),
	   o_Energy_Bin_767      =>   energy_bin_neg_data(766 ),
	   o_Energy_Bin_768      =>   energy_bin_neg_data(767 ),
	   o_Energy_Bin_769      =>   energy_bin_neg_data(768 ),
	   o_Energy_Bin_770      =>   energy_bin_neg_data(769 ),
	   o_Energy_Bin_771      =>   energy_bin_neg_data(770 ),
	   o_Energy_Bin_772      =>   energy_bin_neg_data(771 ),
	   o_Energy_Bin_773      =>   energy_bin_neg_data(772 ),
	   o_Energy_Bin_774      =>   energy_bin_neg_data(773 ),
	   o_Energy_Bin_775      =>   energy_bin_neg_data(774 ),
	   o_Energy_Bin_776      =>   energy_bin_neg_data(775 ),
	   o_Energy_Bin_777      =>   energy_bin_neg_data(776 ),
	   o_Energy_Bin_778      =>   energy_bin_neg_data(777 ),
	   o_Energy_Bin_779      =>   energy_bin_neg_data(778 ),
	   o_Energy_Bin_780      =>   energy_bin_neg_data(779 ),
	   o_Energy_Bin_781      =>   energy_bin_neg_data(780 ),
	   o_Energy_Bin_782      =>   energy_bin_neg_data(781 ),
	   o_Energy_Bin_783      =>   energy_bin_neg_data(782 ),
	   o_Energy_Bin_784      =>   energy_bin_neg_data(783 ),
	   o_Energy_Bin_785      =>   energy_bin_neg_data(784 ),
	   o_Energy_Bin_786      =>   energy_bin_neg_data(785 ),
	   o_Energy_Bin_787      =>   energy_bin_neg_data(786 ),
	   o_Energy_Bin_788      =>   energy_bin_neg_data(787 ),
	   o_Energy_Bin_789      =>   energy_bin_neg_data(788 ),
	   o_Energy_Bin_790      =>   energy_bin_neg_data(789 ),
	   o_Energy_Bin_791      =>   energy_bin_neg_data(790 ),
	   o_Energy_Bin_792      =>   energy_bin_neg_data(791 ),
	   o_Energy_Bin_793      =>   energy_bin_neg_data(792 ),
	   o_Energy_Bin_794      =>   energy_bin_neg_data(793 ),
	   o_Energy_Bin_795      =>   energy_bin_neg_data(794 ),
	   o_Energy_Bin_796      =>   energy_bin_neg_data(795 ),
	   o_Energy_Bin_797      =>   energy_bin_neg_data(796 ),
	   o_Energy_Bin_798      =>   energy_bin_neg_data(797 ),
	   o_Energy_Bin_799      =>   energy_bin_neg_data(798 ),
	   o_Energy_Bin_800      =>   energy_bin_neg_data(799 ),
	   o_Energy_Bin_801      =>   energy_bin_neg_data(800 ),
	   o_Energy_Bin_802      =>   energy_bin_neg_data(801 ),
	   o_Energy_Bin_803      =>   energy_bin_neg_data(802 ),
	   o_Energy_Bin_804      =>   energy_bin_neg_data(803 ),
	   o_Energy_Bin_805      =>   energy_bin_neg_data(804 ),
	   o_Energy_Bin_806      =>   energy_bin_neg_data(805 ),
	   o_Energy_Bin_807      =>   energy_bin_neg_data(806 ),
	   o_Energy_Bin_808      =>   energy_bin_neg_data(807 ),
	   o_Energy_Bin_809      =>   energy_bin_neg_data(808 ),
	   o_Energy_Bin_810      =>   energy_bin_neg_data(809 ),
	   o_Energy_Bin_811      =>   energy_bin_neg_data(810 ),
	   o_Energy_Bin_812      =>   energy_bin_neg_data(811 ),
	   o_Energy_Bin_813      =>   energy_bin_neg_data(812 ),
	   o_Energy_Bin_814      =>   energy_bin_neg_data(813 ),
	   o_Energy_Bin_815      =>   energy_bin_neg_data(814 ),
	   o_Energy_Bin_816      =>   energy_bin_neg_data(815 ),
	   o_Energy_Bin_817      =>   energy_bin_neg_data(816 ),
	   o_Energy_Bin_818      =>   energy_bin_neg_data(817 ),
	   o_Energy_Bin_819      =>   energy_bin_neg_data(818 ),
	   o_Energy_Bin_820      =>   energy_bin_neg_data(819 ),
	   o_Energy_Bin_821      =>   energy_bin_neg_data(820 ),
	   o_Energy_Bin_822      =>   energy_bin_neg_data(821 ),
	   o_Energy_Bin_823      =>   energy_bin_neg_data(822 ),
	   o_Energy_Bin_824      =>   energy_bin_neg_data(823 ),
	   o_Energy_Bin_825      =>   energy_bin_neg_data(824 ),
	   o_Energy_Bin_826      =>   energy_bin_neg_data(825 ),
	   o_Energy_Bin_827      =>   energy_bin_neg_data(826 ),
	   o_Energy_Bin_828      =>   energy_bin_neg_data(827 ),
	   o_Energy_Bin_829      =>   energy_bin_neg_data(828 ),
	   o_Energy_Bin_830      =>   energy_bin_neg_data(829 ),
	   o_Energy_Bin_831      =>   energy_bin_neg_data(830 ),
	   o_Energy_Bin_832      =>   energy_bin_neg_data(831 ),
	   o_Energy_Bin_833      =>   energy_bin_neg_data(832 ),
	   o_Energy_Bin_834      =>   energy_bin_neg_data(833 ),
	   o_Energy_Bin_835      =>   energy_bin_neg_data(834 ),
	   o_Energy_Bin_836      =>   energy_bin_neg_data(835 ),
	   o_Energy_Bin_837      =>   energy_bin_neg_data(836 ),
	   o_Energy_Bin_838      =>   energy_bin_neg_data(837 ),
	   o_Energy_Bin_839      =>   energy_bin_neg_data(838 ),
	   o_Energy_Bin_840      =>   energy_bin_neg_data(839 ),
	   o_Energy_Bin_841      =>   energy_bin_neg_data(840 ),
	   o_Energy_Bin_842      =>   energy_bin_neg_data(841 ),
	   o_Energy_Bin_843      =>   energy_bin_neg_data(842 ),
	   o_Energy_Bin_844      =>   energy_bin_neg_data(843 ),
	   o_Energy_Bin_845      =>   energy_bin_neg_data(844 ),
	   o_Energy_Bin_846      =>   energy_bin_neg_data(845 ),
	   o_Energy_Bin_847      =>   energy_bin_neg_data(846 ),
	   o_Energy_Bin_848      =>   energy_bin_neg_data(847 ),
	   o_Energy_Bin_849      =>   energy_bin_neg_data(848 ),
	   o_Energy_Bin_850      =>   energy_bin_neg_data(849 ),
	   o_Energy_Bin_851      =>   energy_bin_neg_data(850 ),
	   o_Energy_Bin_852      =>   energy_bin_neg_data(851 ),
	   o_Energy_Bin_853      =>   energy_bin_neg_data(852 ),
	   o_Energy_Bin_854      =>   energy_bin_neg_data(853 ),
	   o_Energy_Bin_855      =>   energy_bin_neg_data(854 ),
	   o_Energy_Bin_856      =>   energy_bin_neg_data(855 ),
	   o_Energy_Bin_857      =>   energy_bin_neg_data(856 ),
	   o_Energy_Bin_858      =>   energy_bin_neg_data(857 ),
	   o_Energy_Bin_859      =>   energy_bin_neg_data(858 ),
	   o_Energy_Bin_860      =>   energy_bin_neg_data(859 ),
	   o_Energy_Bin_861      =>   energy_bin_neg_data(860 ),
	   o_Energy_Bin_862      =>   energy_bin_neg_data(861 ),
	   o_Energy_Bin_863      =>   energy_bin_neg_data(862 ),
	   o_Energy_Bin_864      =>   energy_bin_neg_data(863 ),
	   o_Energy_Bin_865      =>   energy_bin_neg_data(864 ),
	   o_Energy_Bin_866      =>   energy_bin_neg_data(865 ),
	   o_Energy_Bin_867      =>   energy_bin_neg_data(866 ),
	   o_Energy_Bin_868      =>   energy_bin_neg_data(867 ),
	   o_Energy_Bin_869      =>   energy_bin_neg_data(868 ),
	   o_Energy_Bin_870      =>   energy_bin_neg_data(869 ),
	   o_Energy_Bin_871      =>   energy_bin_neg_data(870 ),
	   o_Energy_Bin_872      =>   energy_bin_neg_data(871 ),
	   o_Energy_Bin_873      =>   energy_bin_neg_data(872 ),
	   o_Energy_Bin_874      =>   energy_bin_neg_data(873 ),
	   o_Energy_Bin_875      =>   energy_bin_neg_data(874 ),
	   o_Energy_Bin_876      =>   energy_bin_neg_data(875 ),
	   o_Energy_Bin_877      =>   energy_bin_neg_data(876 ),
	   o_Energy_Bin_878      =>   energy_bin_neg_data(877 ),
	   o_Energy_Bin_879      =>   energy_bin_neg_data(878 ),
	   o_Energy_Bin_880      =>   energy_bin_neg_data(879 ),
	   o_Energy_Bin_881      =>   energy_bin_neg_data(880 ),
	   o_Energy_Bin_882      =>   energy_bin_neg_data(881 ),
	   o_Energy_Bin_883      =>   energy_bin_neg_data(882 ),
	   o_Energy_Bin_884      =>   energy_bin_neg_data(883 ),
	   o_Energy_Bin_885      =>   energy_bin_neg_data(884 ),
	   o_Energy_Bin_886      =>   energy_bin_neg_data(885 ),
	   o_Energy_Bin_887      =>   energy_bin_neg_data(886 ),
	   o_Energy_Bin_888      =>   energy_bin_neg_data(887 ),
	   o_Energy_Bin_889      =>   energy_bin_neg_data(888 ),
	   o_Energy_Bin_890      =>   energy_bin_neg_data(889 ),
	   o_Energy_Bin_891      =>   energy_bin_neg_data(890 ),
	   o_Energy_Bin_892      =>   energy_bin_neg_data(891 ),
	   o_Energy_Bin_893      =>   energy_bin_neg_data(892 ),
	   o_Energy_Bin_894      =>   energy_bin_neg_data(893 ),
	   o_Energy_Bin_895      =>   energy_bin_neg_data(894 ),
	   o_Energy_Bin_896      =>   energy_bin_neg_data(895 ),
	   o_Energy_Bin_897      =>   energy_bin_neg_data(896 ),
	   o_Energy_Bin_898      =>   energy_bin_neg_data(897 ),
	   o_Energy_Bin_899      =>   energy_bin_neg_data(898 ),
	   o_Energy_Bin_900      =>   energy_bin_neg_data(899 ),
	   o_Energy_Bin_901      =>   energy_bin_neg_data(900 ),
	   o_Energy_Bin_902      =>   energy_bin_neg_data(901 ),
	   o_Energy_Bin_903      =>   energy_bin_neg_data(902 ),
	   o_Energy_Bin_904      =>   energy_bin_neg_data(903 ),
	   o_Energy_Bin_905      =>   energy_bin_neg_data(904 ),
	   o_Energy_Bin_906      =>   energy_bin_neg_data(905 ),
	   o_Energy_Bin_907      =>   energy_bin_neg_data(906 ),
	   o_Energy_Bin_908      =>   energy_bin_neg_data(907 ),
	   o_Energy_Bin_909      =>   energy_bin_neg_data(908 ),
	   o_Energy_Bin_910      =>   energy_bin_neg_data(909 ),
	   o_Energy_Bin_911      =>   energy_bin_neg_data(910 ),
	   o_Energy_Bin_912      =>   energy_bin_neg_data(911 ),
	   o_Energy_Bin_913      =>   energy_bin_neg_data(912 ),
	   o_Energy_Bin_914      =>   energy_bin_neg_data(913 ),
	   o_Energy_Bin_915      =>   energy_bin_neg_data(914 ),
	   o_Energy_Bin_916      =>   energy_bin_neg_data(915 ),
	   o_Energy_Bin_917      =>   energy_bin_neg_data(916 ),
	   o_Energy_Bin_918      =>   energy_bin_neg_data(917 ),
	   o_Energy_Bin_919      =>   energy_bin_neg_data(918 ),
	   o_Energy_Bin_920      =>   energy_bin_neg_data(919 ),
	   o_Energy_Bin_921      =>   energy_bin_neg_data(920 ),
	   o_Energy_Bin_922      =>   energy_bin_neg_data(921 ),
	   o_Energy_Bin_923      =>   energy_bin_neg_data(922 ),
	   o_Energy_Bin_924      =>   energy_bin_neg_data(923 ),
	   o_Energy_Bin_925      =>   energy_bin_neg_data(924 ),
	   o_Energy_Bin_926      =>   energy_bin_neg_data(925 ),
	   o_Energy_Bin_927      =>   energy_bin_neg_data(926 ),
	   o_Energy_Bin_928      =>   energy_bin_neg_data(927 ),
	   o_Energy_Bin_929      =>   energy_bin_neg_data(928 ),
	   o_Energy_Bin_930      =>   energy_bin_neg_data(929 ),
	   o_Energy_Bin_931      =>   energy_bin_neg_data(930 ),
	   o_Energy_Bin_932      =>   energy_bin_neg_data(931 ),
	   o_Energy_Bin_933      =>   energy_bin_neg_data(932 ),
	   o_Energy_Bin_934      =>   energy_bin_neg_data(933 ),
	   o_Energy_Bin_935      =>   energy_bin_neg_data(934 ),
	   o_Energy_Bin_936      =>   energy_bin_neg_data(935 ),
	   o_Energy_Bin_937      =>   energy_bin_neg_data(936 ),
	   o_Energy_Bin_938      =>   energy_bin_neg_data(937 ),
	   o_Energy_Bin_939      =>   energy_bin_neg_data(938 ),
	   o_Energy_Bin_940      =>   energy_bin_neg_data(939 ),
	   o_Energy_Bin_941      =>   energy_bin_neg_data(940 ),
	   o_Energy_Bin_942      =>   energy_bin_neg_data(941 ),
	   o_Energy_Bin_943      =>   energy_bin_neg_data(942 ),
	   o_Energy_Bin_944      =>   energy_bin_neg_data(943 ),
	   o_Energy_Bin_945      =>   energy_bin_neg_data(944 ),
	   o_Energy_Bin_946      =>   energy_bin_neg_data(945 ),
	   o_Energy_Bin_947      =>   energy_bin_neg_data(946 ),
	   o_Energy_Bin_948      =>   energy_bin_neg_data(947 ),
	   o_Energy_Bin_949      =>   energy_bin_neg_data(948 ),
	   o_Energy_Bin_950      =>   energy_bin_neg_data(949 ),
	   o_Energy_Bin_951      =>   energy_bin_neg_data(950 ),
	   o_Energy_Bin_952      =>   energy_bin_neg_data(951 ),
	   o_Energy_Bin_953      =>   energy_bin_neg_data(952 ),
	   o_Energy_Bin_954      =>   energy_bin_neg_data(953 ),
	   o_Energy_Bin_955      =>   energy_bin_neg_data(954 ),
	   o_Energy_Bin_956      =>   energy_bin_neg_data(955 ),
	   o_Energy_Bin_957      =>   energy_bin_neg_data(956 ),
	   o_Energy_Bin_958      =>   energy_bin_neg_data(957 ),
	   o_Energy_Bin_959      =>   energy_bin_neg_data(958 ),
	   o_Energy_Bin_960      =>   energy_bin_neg_data(959 ),
	   o_Energy_Bin_961      =>   energy_bin_neg_data(960 ),
	   o_Energy_Bin_962      =>   energy_bin_neg_data(961 ),
	   o_Energy_Bin_963      =>   energy_bin_neg_data(962 ),
	   o_Energy_Bin_964      =>   energy_bin_neg_data(963 ),
	   o_Energy_Bin_965      =>   energy_bin_neg_data(964 ),
	   o_Energy_Bin_966      =>   energy_bin_neg_data(965 ),
	   o_Energy_Bin_967      =>   energy_bin_neg_data(966 ),
	   o_Energy_Bin_968      =>   energy_bin_neg_data(967 ),
	   o_Energy_Bin_969      =>   energy_bin_neg_data(968 ),
	   o_Energy_Bin_970      =>   energy_bin_neg_data(969 ),
	   o_Energy_Bin_971      =>   energy_bin_neg_data(970 ),
	   o_Energy_Bin_972      =>   energy_bin_neg_data(971 ),
	   o_Energy_Bin_973      =>   energy_bin_neg_data(972 ),
	   o_Energy_Bin_974      =>   energy_bin_neg_data(973 ),
	   o_Energy_Bin_975      =>   energy_bin_neg_data(974 ),
	   o_Energy_Bin_976      =>   energy_bin_neg_data(975 ),
	   o_Energy_Bin_977      =>   energy_bin_neg_data(976 ),
	   o_Energy_Bin_978      =>   energy_bin_neg_data(977 ),
	   o_Energy_Bin_979      =>   energy_bin_neg_data(978 ),
	   o_Energy_Bin_980      =>   energy_bin_neg_data(979 ),
	   o_Energy_Bin_981      =>   energy_bin_neg_data(980 ),
	   o_Energy_Bin_982      =>   energy_bin_neg_data(981 ),
	   o_Energy_Bin_983      =>   energy_bin_neg_data(982 ),
	   o_Energy_Bin_984      =>   energy_bin_neg_data(983 ),
	   o_Energy_Bin_985      =>   energy_bin_neg_data(984 ),
	   o_Energy_Bin_986      =>   energy_bin_neg_data(985 ),
	   o_Energy_Bin_987      =>   energy_bin_neg_data(986 ),
	   o_Energy_Bin_988      =>   energy_bin_neg_data(987 ),
	   o_Energy_Bin_989      =>   energy_bin_neg_data(988 ),
	   o_Energy_Bin_990      =>   energy_bin_neg_data(989 ),
	   o_Energy_Bin_991      =>   energy_bin_neg_data(990 ),
	   o_Energy_Bin_992      =>   energy_bin_neg_data(991 ),
	   o_Energy_Bin_993      =>   energy_bin_neg_data(992 ),
	   o_Energy_Bin_994      =>   energy_bin_neg_data(993 ),
	   o_Energy_Bin_995      =>   energy_bin_neg_data(994 ),
	   o_Energy_Bin_996      =>   energy_bin_neg_data(995 ),
	   o_Energy_Bin_997      =>   energy_bin_neg_data(996 ),
	   o_Energy_Bin_998      =>   energy_bin_neg_data(997 ),
	   o_Energy_Bin_999      =>   energy_bin_neg_data(998 ),
	   o_Energy_Bin_1000     =>   energy_bin_neg_data(999 ),
	   o_Energy_Bin_1001     =>   energy_bin_neg_data(1000),
	   o_Energy_Bin_1002     =>   energy_bin_neg_data(1001),
	   o_Energy_Bin_1003     =>   energy_bin_neg_data(1002),
	   o_Energy_Bin_1004     =>   energy_bin_neg_data(1003),
	   o_Energy_Bin_1005     =>   energy_bin_neg_data(1004),
	   o_Energy_Bin_1006     =>   energy_bin_neg_data(1005),
	   o_Energy_Bin_1007     =>   energy_bin_neg_data(1006),
	   o_Energy_Bin_1008     =>   energy_bin_neg_data(1007),
	   o_Energy_Bin_1009     =>   energy_bin_neg_data(1008),
	   o_Energy_Bin_1010     =>   energy_bin_neg_data(1009),
	   o_Energy_Bin_1011     =>   energy_bin_neg_data(1010),
	   o_Energy_Bin_1012     =>   energy_bin_neg_data(1011),
	   o_Energy_Bin_1013     =>   energy_bin_neg_data(1012),
	   o_Energy_Bin_1014     =>   energy_bin_neg_data(1013),
	   o_Energy_Bin_1015     =>   energy_bin_neg_data(1014),
	   o_Energy_Bin_1016     =>   energy_bin_neg_data(1015),
	   o_Energy_Bin_1017     =>   energy_bin_neg_data(1016),
	   o_Energy_Bin_1018     =>   energy_bin_neg_data(1017),
	   o_Energy_Bin_1019     =>   energy_bin_neg_data(1018),
	   o_Energy_Bin_1020     =>   energy_bin_neg_data(1019),
	   o_Energy_Bin_1021     =>   energy_bin_neg_data(1020),
	   o_Energy_Bin_1022     =>   energy_bin_neg_data(1021),
	   o_Energy_Bin_1023     =>   energy_bin_neg_data(1022),
	   o_Energy_Bin_1024     =>   energy_bin_neg_data(1023),

       i_PEAK_THD_pos        =>   i_PEAK_THD_pos,
	   i_PEAK_THD            =>   i_PEAK_THD

         );
ReadAdc_inst : TB_ReadAdc
  port map  (
       CLK100       =>    CLK100,
       RST          =>    RST,
       
       ADC_CLK_1    =>    ADC_CLK_1,   
       ADC_CLK_2    =>    ADC_CLK_2,

       ADC_D1     =>   ADC_D1_s   ,
       ADC_DR1    =>   ADC_DR1_s  ,

       ADC_D2     =>   ADC_D2_s   ,
       ADC_DR2    =>   ADC_DR2_s  ,
       
       i_DR1_EN     =>   i_DR1_EN,
       i_DR2_EN     =>   i_DR2_EN,
       
       DATA1      =>   DATA1    ,
       DATARDY1   =>   DATARDY1 ,  
       DATA2      =>   DATA2    ,
       DATARDY2   =>   DATARDY2 ,
	   
	   i_stop_req =>   i_stop_req
        );
        
--adc raw data fifos control ***********************************************************************************************************************************************************************************
adc_fifo_ctrl_tlm_1: process (CLK100, RST)
begin
  if RST = '1' then
        wr_en_adc_fifo_1  <= '0';
        energy_bin_cnt_1  <= 0;
  elsif rising_edge(CLK100) then
        if( mtime_over = '1' and adc_fifo_full_1 = '0' and energy_bin_cnt_1 < 1024) then
            energy_bin_cnt_1 <= energy_bin_cnt_1 + 1;
            wr_en_adc_fifo_1  <= '1';
            adc_fifo_data_in_1 <= energy_bin_pos_data(energy_bin_cnt_1);
        else
            wr_en_adc_fifo_1  <= '0';
        end if;
    
  end if;
end process;

adc_fifo_ctrl_tlm_2: process (CLK100, RST)
begin
  if RST = '1' then
        wr_en_adc_fifo_2  <= '0';
        energy_bin_cnt_2  <= 0;
  elsif rising_edge(CLK100) then
        if( mtime_over = '1' and adc_fifo_full_2 = '0' and energy_bin_cnt_2 < 1024) then
            energy_bin_cnt_2 <= energy_bin_cnt_2 + 1;
            wr_en_adc_fifo_2  <= '1';
            adc_fifo_data_in_2 <= energy_bin_neg_data(energy_bin_cnt_2);
        else
            wr_en_adc_fifo_2  <= '0';
        end if;
    
  end if;
end process;

-- peak fifos ************************************************************************************************************************************************************************************************

peak_fifo_ctrl_tlm_1: process (CLK100, RST)
begin
  if RST = '1' then
        wr_en_peak_fifo_1  <= '0';
        peak_fifo_wr_cnt_1 <= (others => '0');
  elsif rising_edge(CLK100) then
        if( PEAK_FL_C1_s = '1' and peak_fifo_full_1 = '0' and peak_fifo_wr_cnt_1 < 2001) then
            peak_fifo_wr_cnt_1 <= peak_fifo_wr_cnt_1 + '1';
            wr_en_peak_fifo_1  <= '1';
            peak_fifo_data_in_1 <= PEAK_C1_s;
        else
            wr_en_peak_fifo_1  <= '0';
        end if;
    
  end if;
end process;

peak_fifo_ctrl_tlm_2: process (CLK100, RST)
begin
  if RST = '1' then
        wr_en_peak_fifo_2  <= '0';
        peak_fifo_wr_cnt_2 <= (others => '0');
  elsif rising_edge(CLK100) then
        if( PEAK_FL_C1_s_pos = '1' and peak_fifo_full_2 = '0' and peak_fifo_wr_cnt_2 < 2001) then
            peak_fifo_wr_cnt_2 <= peak_fifo_wr_cnt_2 + '1';
            wr_en_peak_fifo_2  <= '1';
            peak_fifo_data_in_2 <= PEAK_C1_s_pos;
        else
            wr_en_peak_fifo_2  <= '0';
        end if;
    
  end if;
end process;
          
end architecture DataCtrl_RTL;
--============================================================================
-- Architecture definition section end - RTL
--****************************************************************************


--****************************************************************************
-- Module trailer section starts
--============================================================================
--
--
--
--
--
--============================================================================
-- Module trailer section ends
--****************************************************************************


