-- Copyright reserved University of Alberta
--Author: Bo Yu
--+----------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.numeric_STD.all;


entity PeakDetector is
  --+----------
  -- Generic declarations
  --+----------
  generic(                        
        DataVecSize_g  		      :integer := 56;
        WdVecSize_g    		      :integer := 16;
        ByteSize_g     		      :integer := 8;
        NibbleSize_g   		      :integer := 4; 

		s_E1_C1_L        	 	  :std_logic_vector(11 downto 0) := x"000"; 
		s_E1_C1_H        	 	  :std_logic_vector(11 downto 0) := x"002"; 
		s_E2_C1_H        	 	  :std_logic_vector(11 downto 0) := x"004"; 
		s_E3_C1_H        	 	  :std_logic_vector(11 downto 0) := x"006"; 
		s_E4_C1_H        	 	  :std_logic_vector(11 downto 0) := x"008"; 
		s_E5_C1_H        	 	  :std_logic_vector(11 downto 0) := x"00A"; 
		s_E6_C1_H        	 	  :std_logic_vector(11 downto 0) := x"00C"; 
		s_E7_C1_H        	 	  :std_logic_vector(11 downto 0) := x"00E"; 
		s_E8_C1_H        	 	  :std_logic_vector(11 downto 0) := x"010"; 
		s_E9_C1_H        	 	  :std_logic_vector(11 downto 0) := x"012"; 
		s_E10_C1_H       	 	  :std_logic_vector(11 downto 0) := x"014"; 
		s_E11_C1_H				  :std_logic_vector(11 downto 0) := x"016"; 
		s_E12_C1_H				  :std_logic_vector(11 downto 0) := x"018"; 
		s_E13_C1_H				  :std_logic_vector(11 downto 0) := x"01A"; 
		s_E14_C1_H				  :std_logic_vector(11 downto 0) := x"01C"; 
		s_E15_C1_H				  :std_logic_vector(11 downto 0) := x"01E"; 
		s_E16_C1_H				  :std_logic_vector(11 downto 0) := x"020"; 
		s_E17_C1_H				  :std_logic_vector(11 downto 0) := x"022"; 
		s_E18_C1_H				  :std_logic_vector(11 downto 0) := x"024"; 
		s_E19_C1_H				  :std_logic_vector(11 downto 0) := x"026"; 
		s_E20_C1_H				  :std_logic_vector(11 downto 0) := x"028"; 
		s_E21_C1_H				  :std_logic_vector(11 downto 0) := x"02A"; 
		s_E22_C1_H				  :std_logic_vector(11 downto 0) := x"02C"; 
		s_E23_C1_H				  :std_logic_vector(11 downto 0) := x"02E"; 
		s_E24_C1_H				  :std_logic_vector(11 downto 0) := x"030"; 
		s_E25_C1_H				  :std_logic_vector(11 downto 0) := x"032"; 
		s_E26_C1_H				  :std_logic_vector(11 downto 0) := x"034"; 
		s_E27_C1_H				  :std_logic_vector(11 downto 0) := x"036"; 
		s_E28_C1_H				  :std_logic_vector(11 downto 0) := x"038"; 
		s_E29_C1_H				  :std_logic_vector(11 downto 0) := x"03A"; 
		s_E30_C1_H				  :std_logic_vector(11 downto 0) := x"03C"; 
		s_E31_C1_H				  :std_logic_vector(11 downto 0) := x"03E"; 
		s_E32_C1_H				  :std_logic_vector(11 downto 0) := x"040"; 
		s_E33_C1_H				  :std_logic_vector(11 downto 0) := x"042"; 
		s_E34_C1_H				  :std_logic_vector(11 downto 0) := x"044"; 
		s_E35_C1_H				  :std_logic_vector(11 downto 0) := x"046"; 
		s_E36_C1_H				  :std_logic_vector(11 downto 0) := x"048"; 
		s_E37_C1_H				  :std_logic_vector(11 downto 0) := x"04A"; 
		s_E38_C1_H				  :std_logic_vector(11 downto 0) := x"04C"; 
		s_E39_C1_H				  :std_logic_vector(11 downto 0) := x"04E"; 
		s_E40_C1_H				  :std_logic_vector(11 downto 0) := x"050"; 
		s_E41_C1_H				  :std_logic_vector(11 downto 0) := x"052"; 
		s_E42_C1_H				  :std_logic_vector(11 downto 0) := x"054"; 
		s_E43_C1_H				  :std_logic_vector(11 downto 0) := x"056"; 
		s_E44_C1_H				  :std_logic_vector(11 downto 0) := x"058"; 
		s_E45_C1_H				  :std_logic_vector(11 downto 0) := x"05A"; 
		s_E46_C1_H				  :std_logic_vector(11 downto 0) := x"05C"; 
		s_E47_C1_H				  :std_logic_vector(11 downto 0) := x"05E"; 
		s_E48_C1_H				  :std_logic_vector(11 downto 0) := x"060"; 
		s_E49_C1_H				  :std_logic_vector(11 downto 0) := x"062"; 
		s_E50_C1_H				  :std_logic_vector(11 downto 0) := x"064"; 
		s_E51_C1_H				  :std_logic_vector(11 downto 0) := x"066"; 
		s_E52_C1_H				  :std_logic_vector(11 downto 0) := x"068"; 
		s_E53_C1_H				  :std_logic_vector(11 downto 0) := x"06A"; 
		s_E54_C1_H				  :std_logic_vector(11 downto 0) := x"06C"; 
		s_E55_C1_H				  :std_logic_vector(11 downto 0) := x"06E"; 
		s_E56_C1_H				  :std_logic_vector(11 downto 0) := x"070"; 
		s_E57_C1_H				  :std_logic_vector(11 downto 0) := x"072"; 
		s_E58_C1_H				  :std_logic_vector(11 downto 0) := x"074"; 
		s_E59_C1_H				  :std_logic_vector(11 downto 0) := x"076"; 
		s_E60_C1_H				  :std_logic_vector(11 downto 0) := x"078"; 
		s_E61_C1_H				  :std_logic_vector(11 downto 0) := x"07A"; 
		s_E62_C1_H				  :std_logic_vector(11 downto 0) := x"07C"; 
		s_E63_C1_H				  :std_logic_vector(11 downto 0) := x"07E"; 
		s_E64_C1_H				  :std_logic_vector(11 downto 0) := x"080"; 
		s_E65_C1_H				  :std_logic_vector(11 downto 0) := x"082"; 
		s_E66_C1_H				  :std_logic_vector(11 downto 0) := x"084"; 
		s_E67_C1_H				  :std_logic_vector(11 downto 0) := x"086"; 
		s_E68_C1_H				  :std_logic_vector(11 downto 0) := x"088"; 
		s_E69_C1_H				  :std_logic_vector(11 downto 0) := x"08A"; 
		s_E70_C1_H				  :std_logic_vector(11 downto 0) := x"08C"; 
		s_E71_C1_H				  :std_logic_vector(11 downto 0) := x"08E"; 
		s_E72_C1_H				  :std_logic_vector(11 downto 0) := x"090"; 
		s_E73_C1_H				  :std_logic_vector(11 downto 0) := x"092"; 
		s_E74_C1_H				  :std_logic_vector(11 downto 0) := x"094"; 
		s_E75_C1_H				  :std_logic_vector(11 downto 0) := x"096"; 
		s_E76_C1_H				  :std_logic_vector(11 downto 0) := x"098"; 
		s_E77_C1_H				  :std_logic_vector(11 downto 0) := x"09A"; 
		s_E78_C1_H				  :std_logic_vector(11 downto 0) := x"09C"; 
		s_E79_C1_H				  :std_logic_vector(11 downto 0) := x"09E"; 
		s_E80_C1_H				  :std_logic_vector(11 downto 0) := x"0A0"; 
		s_E81_C1_H				  :std_logic_vector(11 downto 0) := x"0A2"; 
		s_E82_C1_H				  :std_logic_vector(11 downto 0) := x"0A4"; 
		s_E83_C1_H				  :std_logic_vector(11 downto 0) := x"0A6"; 
		s_E84_C1_H				  :std_logic_vector(11 downto 0) := x"0A8"; 
		s_E85_C1_H				  :std_logic_vector(11 downto 0) := x"0AA"; 
		s_E86_C1_H				  :std_logic_vector(11 downto 0) := x"0AC"; 
		s_E87_C1_H				  :std_logic_vector(11 downto 0) := x"0AE"; 
		s_E88_C1_H				  :std_logic_vector(11 downto 0) := x"0B0"; 
		s_E89_C1_H				  :std_logic_vector(11 downto 0) := x"0B2"; 
		s_E90_C1_H				  :std_logic_vector(11 downto 0) := x"0B4"; 
		s_E91_C1_H				  :std_logic_vector(11 downto 0) := x"0B6"; 
		s_E92_C1_H				  :std_logic_vector(11 downto 0) := x"0B8"; 
		s_E93_C1_H				  :std_logic_vector(11 downto 0) := x"0BA"; 
		s_E94_C1_H				  :std_logic_vector(11 downto 0) := x"0BC"; 
		s_E95_C1_H				  :std_logic_vector(11 downto 0) := x"0BE"; 
		s_E96_C1_H				  :std_logic_vector(11 downto 0) := x"0C0"; 
		s_E97_C1_H				  :std_logic_vector(11 downto 0) := x"0C2"; 
		s_E98_C1_H				  :std_logic_vector(11 downto 0) := x"0C4"; 
		s_E99_C1_H				  :std_logic_vector(11 downto 0) := x"0C6"; 
		s_E100_C1_H				  :std_logic_vector(11 downto 0) := x"0C8"; 
		s_E101_C1_H				  :std_logic_vector(11 downto 0) := x"0CA"; 
		s_E102_C1_H				  :std_logic_vector(11 downto 0) := x"0CC"; 
		s_E103_C1_H				  :std_logic_vector(11 downto 0) := x"0CE"; 
		s_E104_C1_H				  :std_logic_vector(11 downto 0) := x"0D0"; 
		s_E105_C1_H				  :std_logic_vector(11 downto 0) := x"0D2"; 
		s_E106_C1_H				  :std_logic_vector(11 downto 0) := x"0D4"; 
		s_E107_C1_H				  :std_logic_vector(11 downto 0) := x"0D6"; 
		s_E108_C1_H				  :std_logic_vector(11 downto 0) := x"0D8"; 
		s_E109_C1_H				  :std_logic_vector(11 downto 0) := x"0DA"; 
		s_E110_C1_H				  :std_logic_vector(11 downto 0) := x"0DC"; 
		s_E111_C1_H				  :std_logic_vector(11 downto 0) := x"0DE"; 
		s_E112_C1_H				  :std_logic_vector(11 downto 0) := x"0E0"; 
		s_E113_C1_H				  :std_logic_vector(11 downto 0) := x"0E2"; 
		s_E114_C1_H				  :std_logic_vector(11 downto 0) := x"0E4"; 
		s_E115_C1_H				  :std_logic_vector(11 downto 0) := x"0E6"; 
		s_E116_C1_H				  :std_logic_vector(11 downto 0) := x"0E8"; 
		s_E117_C1_H				  :std_logic_vector(11 downto 0) := x"0EA"; 
		s_E118_C1_H				  :std_logic_vector(11 downto 0) := x"0EC"; 
		s_E119_C1_H				  :std_logic_vector(11 downto 0) := x"0EE"; 
		s_E120_C1_H				  :std_logic_vector(11 downto 0) := x"0F0"; 
		s_E121_C1_H				  :std_logic_vector(11 downto 0) := x"0F2"; 
		s_E122_C1_H				  :std_logic_vector(11 downto 0) := x"0F4"; 
		s_E123_C1_H				  :std_logic_vector(11 downto 0) := x"0F6"; 
		s_E124_C1_H				  :std_logic_vector(11 downto 0) := x"0F8"; 
		s_E125_C1_H				  :std_logic_vector(11 downto 0) := x"0FA"; 
		s_E126_C1_H				  :std_logic_vector(11 downto 0) := x"0FC"; 
		s_E127_C1_H				  :std_logic_vector(11 downto 0) := x"0FE"; 
		s_E128_C1_H				  :std_logic_vector(11 downto 0) := x"100"; 
		s_E129_C1_H				  :std_logic_vector(11 downto 0) := x"102"; 
		s_E130_C1_H				  :std_logic_vector(11 downto 0) := x"104"; 
		s_E131_C1_H				  :std_logic_vector(11 downto 0) := x"106"; 
		s_E132_C1_H				  :std_logic_vector(11 downto 0) := x"108"; 
		s_E133_C1_H				  :std_logic_vector(11 downto 0) := x"10A"; 
		s_E134_C1_H				  :std_logic_vector(11 downto 0) := x"10C"; 
		s_E135_C1_H				  :std_logic_vector(11 downto 0) := x"10E"; 
		s_E136_C1_H				  :std_logic_vector(11 downto 0) := x"110"; 
		s_E137_C1_H				  :std_logic_vector(11 downto 0) := x"112"; 
		s_E138_C1_H				  :std_logic_vector(11 downto 0) := x"114"; 
		s_E139_C1_H				  :std_logic_vector(11 downto 0) := x"116"; 
		s_E140_C1_H				  :std_logic_vector(11 downto 0) := x"118"; 
		s_E141_C1_H				  :std_logic_vector(11 downto 0) := x"11A"; 
		s_E142_C1_H				  :std_logic_vector(11 downto 0) := x"11C"; 
		s_E143_C1_H				  :std_logic_vector(11 downto 0) := x"11E"; 
		s_E144_C1_H				  :std_logic_vector(11 downto 0) := x"120"; 
		s_E145_C1_H				  :std_logic_vector(11 downto 0) := x"122"; 
		s_E146_C1_H				  :std_logic_vector(11 downto 0) := x"124"; 
		s_E147_C1_H				  :std_logic_vector(11 downto 0) := x"126"; 
		s_E148_C1_H				  :std_logic_vector(11 downto 0) := x"128"; 
		s_E149_C1_H				  :std_logic_vector(11 downto 0) := x"12A"; 
		s_E150_C1_H				  :std_logic_vector(11 downto 0) := x"12C"; 
		s_E151_C1_H				  :std_logic_vector(11 downto 0) := x"12E"; 
		s_E152_C1_H				  :std_logic_vector(11 downto 0) := x"130"; 
		s_E153_C1_H				  :std_logic_vector(11 downto 0) := x"132"; 
		s_E154_C1_H				  :std_logic_vector(11 downto 0) := x"134"; 
		s_E155_C1_H				  :std_logic_vector(11 downto 0) := x"136"; 
		s_E156_C1_H				  :std_logic_vector(11 downto 0) := x"138"; 
		s_E157_C1_H				  :std_logic_vector(11 downto 0) := x"13A"; 
		s_E158_C1_H				  :std_logic_vector(11 downto 0) := x"13C"; 
		s_E159_C1_H				  :std_logic_vector(11 downto 0) := x"13E"; 
		s_E160_C1_H				  :std_logic_vector(11 downto 0) := x"140"; 
		s_E161_C1_H				  :std_logic_vector(11 downto 0) := x"142"; 
		s_E162_C1_H				  :std_logic_vector(11 downto 0) := x"144"; 
		s_E163_C1_H				  :std_logic_vector(11 downto 0) := x"146"; 
		s_E164_C1_H				  :std_logic_vector(11 downto 0) := x"148"; 
		s_E165_C1_H				  :std_logic_vector(11 downto 0) := x"14A"; 
		s_E166_C1_H				  :std_logic_vector(11 downto 0) := x"14C"; 
		s_E167_C1_H				  :std_logic_vector(11 downto 0) := x"14E"; 
		s_E168_C1_H				  :std_logic_vector(11 downto 0) := x"150"; 
		s_E169_C1_H				  :std_logic_vector(11 downto 0) := x"152"; 
		s_E170_C1_H				  :std_logic_vector(11 downto 0) := x"154"; 
		s_E171_C1_H				  :std_logic_vector(11 downto 0) := x"156"; 
		s_E172_C1_H				  :std_logic_vector(11 downto 0) := x"158"; 
		s_E173_C1_H				  :std_logic_vector(11 downto 0) := x"15A"; 
		s_E174_C1_H				  :std_logic_vector(11 downto 0) := x"15C"; 
		s_E175_C1_H				  :std_logic_vector(11 downto 0) := x"15E"; 
		s_E176_C1_H				  :std_logic_vector(11 downto 0) := x"160"; 
		s_E177_C1_H				  :std_logic_vector(11 downto 0) := x"162"; 
		s_E178_C1_H				  :std_logic_vector(11 downto 0) := x"164"; 
		s_E179_C1_H				  :std_logic_vector(11 downto 0) := x"166"; 
		s_E180_C1_H				  :std_logic_vector(11 downto 0) := x"168"; 
		s_E181_C1_H				  :std_logic_vector(11 downto 0) := x"16A"; 
		s_E182_C1_H				  :std_logic_vector(11 downto 0) := x"16C"; 
		s_E183_C1_H				  :std_logic_vector(11 downto 0) := x"16E"; 
		s_E184_C1_H				  :std_logic_vector(11 downto 0) := x"170"; 
		s_E185_C1_H				  :std_logic_vector(11 downto 0) := x"172"; 
		s_E186_C1_H				  :std_logic_vector(11 downto 0) := x"174"; 
		s_E187_C1_H				  :std_logic_vector(11 downto 0) := x"176"; 
		s_E188_C1_H				  :std_logic_vector(11 downto 0) := x"178"; 
		s_E189_C1_H				  :std_logic_vector(11 downto 0) := x"17A"; 
		s_E190_C1_H				  :std_logic_vector(11 downto 0) := x"17C"; 
		s_E191_C1_H				  :std_logic_vector(11 downto 0) := x"17E"; 
		s_E192_C1_H				  :std_logic_vector(11 downto 0) := x"180"; 
		s_E193_C1_H				  :std_logic_vector(11 downto 0) := x"182"; 
		s_E194_C1_H				  :std_logic_vector(11 downto 0) := x"184"; 
		s_E195_C1_H				  :std_logic_vector(11 downto 0) := x"186"; 
		s_E196_C1_H				  :std_logic_vector(11 downto 0) := x"188"; 
		s_E197_C1_H				  :std_logic_vector(11 downto 0) := x"18A"; 
		s_E198_C1_H				  :std_logic_vector(11 downto 0) := x"18C"; 
		s_E199_C1_H				  :std_logic_vector(11 downto 0) := x"18E"; 
		s_E200_C1_H				  :std_logic_vector(11 downto 0) := x"190"; 
		s_E201_C1_H				  :std_logic_vector(11 downto 0) := x"192"; 
		s_E202_C1_H				  :std_logic_vector(11 downto 0) := x"194"; 
		s_E203_C1_H				  :std_logic_vector(11 downto 0) := x"196"; 
		s_E204_C1_H				  :std_logic_vector(11 downto 0) := x"198"; 
		s_E205_C1_H				  :std_logic_vector(11 downto 0) := x"19A"; 
		s_E206_C1_H				  :std_logic_vector(11 downto 0) := x"19C"; 
		s_E207_C1_H				  :std_logic_vector(11 downto 0) := x"19E"; 
		s_E208_C1_H				  :std_logic_vector(11 downto 0) := x"1A0"; 
		s_E209_C1_H				  :std_logic_vector(11 downto 0) := x"1A2"; 
		s_E210_C1_H				  :std_logic_vector(11 downto 0) := x"1A4"; 
		s_E211_C1_H				  :std_logic_vector(11 downto 0) := x"1A6"; 
		s_E212_C1_H				  :std_logic_vector(11 downto 0) := x"1A8"; 
		s_E213_C1_H				  :std_logic_vector(11 downto 0) := x"1AA"; 
		s_E214_C1_H				  :std_logic_vector(11 downto 0) := x"1AC"; 
		s_E215_C1_H				  :std_logic_vector(11 downto 0) := x"1AE"; 
		s_E216_C1_H				  :std_logic_vector(11 downto 0) := x"1B0"; 
		s_E217_C1_H				  :std_logic_vector(11 downto 0) := x"1B2"; 
		s_E218_C1_H				  :std_logic_vector(11 downto 0) := x"1B4"; 
		s_E219_C1_H				  :std_logic_vector(11 downto 0) := x"1B6"; 
		s_E220_C1_H				  :std_logic_vector(11 downto 0) := x"1B8"; 
		s_E221_C1_H				  :std_logic_vector(11 downto 0) := x"1BA"; 
		s_E222_C1_H				  :std_logic_vector(11 downto 0) := x"1BC"; 
		s_E223_C1_H				  :std_logic_vector(11 downto 0) := x"1BE"; 
		s_E224_C1_H				  :std_logic_vector(11 downto 0) := x"1C0"; 
		s_E225_C1_H				  :std_logic_vector(11 downto 0) := x"1C2"; 
		s_E226_C1_H				  :std_logic_vector(11 downto 0) := x"1C4"; 
		s_E227_C1_H				  :std_logic_vector(11 downto 0) := x"1C6"; 
		s_E228_C1_H				  :std_logic_vector(11 downto 0) := x"1C8"; 
		s_E229_C1_H				  :std_logic_vector(11 downto 0) := x"1CA"; 
		s_E230_C1_H				  :std_logic_vector(11 downto 0) := x"1CC"; 
		s_E231_C1_H				  :std_logic_vector(11 downto 0) := x"1CE"; 
		s_E232_C1_H				  :std_logic_vector(11 downto 0) := x"1D0"; 
		s_E233_C1_H				  :std_logic_vector(11 downto 0) := x"1D2"; 
		s_E234_C1_H				  :std_logic_vector(11 downto 0) := x"1D4"; 
		s_E235_C1_H				  :std_logic_vector(11 downto 0) := x"1D6"; 
		s_E236_C1_H				  :std_logic_vector(11 downto 0) := x"1D8"; 
		s_E237_C1_H				  :std_logic_vector(11 downto 0) := x"1DA"; 
		s_E238_C1_H				  :std_logic_vector(11 downto 0) := x"1DC"; 
		s_E239_C1_H				  :std_logic_vector(11 downto 0) := x"1DE"; 
		s_E240_C1_H				  :std_logic_vector(11 downto 0) := x"1E0"; 
		s_E241_C1_H				  :std_logic_vector(11 downto 0) := x"1E2"; 
		s_E242_C1_H				  :std_logic_vector(11 downto 0) := x"1E4"; 
		s_E243_C1_H				  :std_logic_vector(11 downto 0) := x"1E6"; 
		s_E244_C1_H				  :std_logic_vector(11 downto 0) := x"1E8"; 
		s_E245_C1_H				  :std_logic_vector(11 downto 0) := x"1EA"; 
		s_E246_C1_H				  :std_logic_vector(11 downto 0) := x"1EC"; 
		s_E247_C1_H				  :std_logic_vector(11 downto 0) := x"1EE"; 
		s_E248_C1_H				  :std_logic_vector(11 downto 0) := x"1F0"; 
		s_E249_C1_H				  :std_logic_vector(11 downto 0) := x"1F2"; 
		s_E250_C1_H				  :std_logic_vector(11 downto 0) := x"1F4"; 
		s_E251_C1_H				  :std_logic_vector(11 downto 0) := x"1F6"; 
		s_E252_C1_H				  :std_logic_vector(11 downto 0) := x"1F8"; 
		s_E253_C1_H				  :std_logic_vector(11 downto 0) := x"1FA"; 
		s_E254_C1_H				  :std_logic_vector(11 downto 0) := x"1FC"; 
		s_E255_C1_H				  :std_logic_vector(11 downto 0) := x"1FE"; 
		s_E256_C1_H				  :std_logic_vector(11 downto 0) := x"200"; 
		s_E257_C1_H				  :std_logic_vector(11 downto 0) := x"202"; 
		s_E258_C1_H				  :std_logic_vector(11 downto 0) := x"204"; 
		s_E259_C1_H				  :std_logic_vector(11 downto 0) := x"206"; 
		s_E260_C1_H				  :std_logic_vector(11 downto 0) := x"208"; 
		s_E261_C1_H				  :std_logic_vector(11 downto 0) := x"20A"; 
		s_E262_C1_H				  :std_logic_vector(11 downto 0) := x"20C"; 
		s_E263_C1_H				  :std_logic_vector(11 downto 0) := x"20E"; 
		s_E264_C1_H				  :std_logic_vector(11 downto 0) := x"210"; 
		s_E265_C1_H				  :std_logic_vector(11 downto 0) := x"212"; 
		s_E266_C1_H				  :std_logic_vector(11 downto 0) := x"214"; 
		s_E267_C1_H				  :std_logic_vector(11 downto 0) := x"216"; 
		s_E268_C1_H				  :std_logic_vector(11 downto 0) := x"218"; 
		s_E269_C1_H				  :std_logic_vector(11 downto 0) := x"21A"; 
		s_E270_C1_H				  :std_logic_vector(11 downto 0) := x"21C"; 
		s_E271_C1_H				  :std_logic_vector(11 downto 0) := x"21E"; 
		s_E272_C1_H				  :std_logic_vector(11 downto 0) := x"220"; 
		s_E273_C1_H				  :std_logic_vector(11 downto 0) := x"222"; 
		s_E274_C1_H				  :std_logic_vector(11 downto 0) := x"224"; 
		s_E275_C1_H				  :std_logic_vector(11 downto 0) := x"226"; 
		s_E276_C1_H				  :std_logic_vector(11 downto 0) := x"228"; 
		s_E277_C1_H				  :std_logic_vector(11 downto 0) := x"22A"; 
		s_E278_C1_H				  :std_logic_vector(11 downto 0) := x"22C"; 
		s_E279_C1_H				  :std_logic_vector(11 downto 0) := x"22E"; 
		s_E280_C1_H				  :std_logic_vector(11 downto 0) := x"230"; 
		s_E281_C1_H				  :std_logic_vector(11 downto 0) := x"232"; 
		s_E282_C1_H				  :std_logic_vector(11 downto 0) := x"234"; 
		s_E283_C1_H				  :std_logic_vector(11 downto 0) := x"236"; 
		s_E284_C1_H				  :std_logic_vector(11 downto 0) := x"238"; 
		s_E285_C1_H				  :std_logic_vector(11 downto 0) := x"23A"; 
		s_E286_C1_H				  :std_logic_vector(11 downto 0) := x"23C"; 
		s_E287_C1_H				  :std_logic_vector(11 downto 0) := x"23E"; 
		s_E288_C1_H				  :std_logic_vector(11 downto 0) := x"240"; 
		s_E289_C1_H				  :std_logic_vector(11 downto 0) := x"242"; 
		s_E290_C1_H				  :std_logic_vector(11 downto 0) := x"244"; 
		s_E291_C1_H				  :std_logic_vector(11 downto 0) := x"246"; 
		s_E292_C1_H				  :std_logic_vector(11 downto 0) := x"248"; 
		s_E293_C1_H				  :std_logic_vector(11 downto 0) := x"24A"; 
		s_E294_C1_H				  :std_logic_vector(11 downto 0) := x"24C"; 
		s_E295_C1_H				  :std_logic_vector(11 downto 0) := x"24E"; 
		s_E296_C1_H				  :std_logic_vector(11 downto 0) := x"250"; 
		s_E297_C1_H				  :std_logic_vector(11 downto 0) := x"252"; 
		s_E298_C1_H				  :std_logic_vector(11 downto 0) := x"254"; 
		s_E299_C1_H				  :std_logic_vector(11 downto 0) := x"256"; 
		s_E300_C1_H				  :std_logic_vector(11 downto 0) := x"258"; 
		s_E301_C1_H				  :std_logic_vector(11 downto 0) := x"25A"; 
		s_E302_C1_H				  :std_logic_vector(11 downto 0) := x"25C"; 
		s_E303_C1_H				  :std_logic_vector(11 downto 0) := x"25E"; 
		s_E304_C1_H				  :std_logic_vector(11 downto 0) := x"260"; 
		s_E305_C1_H				  :std_logic_vector(11 downto 0) := x"262"; 
		s_E306_C1_H				  :std_logic_vector(11 downto 0) := x"264"; 
		s_E307_C1_H				  :std_logic_vector(11 downto 0) := x"266"; 
		s_E308_C1_H				  :std_logic_vector(11 downto 0) := x"268"; 
		s_E309_C1_H				  :std_logic_vector(11 downto 0) := x"26A"; 
		s_E310_C1_H				  :std_logic_vector(11 downto 0) := x"26C"; 
		s_E311_C1_H				  :std_logic_vector(11 downto 0) := x"26E"; 
		s_E312_C1_H				  :std_logic_vector(11 downto 0) := x"270"; 
		s_E313_C1_H				  :std_logic_vector(11 downto 0) := x"272"; 
		s_E314_C1_H				  :std_logic_vector(11 downto 0) := x"274"; 
		s_E315_C1_H				  :std_logic_vector(11 downto 0) := x"276"; 
		s_E316_C1_H				  :std_logic_vector(11 downto 0) := x"278"; 
		s_E317_C1_H				  :std_logic_vector(11 downto 0) := x"27A"; 
		s_E318_C1_H				  :std_logic_vector(11 downto 0) := x"27C"; 
		s_E319_C1_H				  :std_logic_vector(11 downto 0) := x"27E"; 
		s_E320_C1_H				  :std_logic_vector(11 downto 0) := x"280"; 
		s_E321_C1_H				  :std_logic_vector(11 downto 0) := x"282"; 
		s_E322_C1_H				  :std_logic_vector(11 downto 0) := x"284"; 
		s_E323_C1_H				  :std_logic_vector(11 downto 0) := x"286"; 
		s_E324_C1_H				  :std_logic_vector(11 downto 0) := x"288"; 
		s_E325_C1_H				  :std_logic_vector(11 downto 0) := x"28A"; 
		s_E326_C1_H				  :std_logic_vector(11 downto 0) := x"28C"; 
		s_E327_C1_H				  :std_logic_vector(11 downto 0) := x"28E"; 
		s_E328_C1_H				  :std_logic_vector(11 downto 0) := x"290"; 
		s_E329_C1_H				  :std_logic_vector(11 downto 0) := x"292"; 
		s_E330_C1_H				  :std_logic_vector(11 downto 0) := x"294"; 
		s_E331_C1_H				  :std_logic_vector(11 downto 0) := x"296"; 
		s_E332_C1_H				  :std_logic_vector(11 downto 0) := x"298"; 
		s_E333_C1_H				  :std_logic_vector(11 downto 0) := x"29A"; 
		s_E334_C1_H				  :std_logic_vector(11 downto 0) := x"29C"; 
		s_E335_C1_H				  :std_logic_vector(11 downto 0) := x"29E"; 
		s_E336_C1_H				  :std_logic_vector(11 downto 0) := x"2A0"; 
		s_E337_C1_H				  :std_logic_vector(11 downto 0) := x"2A2"; 
		s_E338_C1_H				  :std_logic_vector(11 downto 0) := x"2A4"; 
		s_E339_C1_H				  :std_logic_vector(11 downto 0) := x"2A6"; 
		s_E340_C1_H				  :std_logic_vector(11 downto 0) := x"2A8"; 
		s_E341_C1_H				  :std_logic_vector(11 downto 0) := x"2AA"; 
		s_E342_C1_H				  :std_logic_vector(11 downto 0) := x"2AC"; 
		s_E343_C1_H				  :std_logic_vector(11 downto 0) := x"2AE"; 
		s_E344_C1_H				  :std_logic_vector(11 downto 0) := x"2B0"; 
		s_E345_C1_H				  :std_logic_vector(11 downto 0) := x"2B2"; 
		s_E346_C1_H				  :std_logic_vector(11 downto 0) := x"2B4"; 
		s_E347_C1_H				  :std_logic_vector(11 downto 0) := x"2B6"; 
		s_E348_C1_H				  :std_logic_vector(11 downto 0) := x"2B8"; 
		s_E349_C1_H				  :std_logic_vector(11 downto 0) := x"2BA"; 
		s_E350_C1_H				  :std_logic_vector(11 downto 0) := x"2BC"; 
		s_E351_C1_H				  :std_logic_vector(11 downto 0) := x"2BE"; 
		s_E352_C1_H				  :std_logic_vector(11 downto 0) := x"2C0"; 
		s_E353_C1_H				  :std_logic_vector(11 downto 0) := x"2C2"; 
		s_E354_C1_H				  :std_logic_vector(11 downto 0) := x"2C4"; 
		s_E355_C1_H				  :std_logic_vector(11 downto 0) := x"2C6"; 
		s_E356_C1_H				  :std_logic_vector(11 downto 0) := x"2C8"; 
		s_E357_C1_H				  :std_logic_vector(11 downto 0) := x"2CA"; 
		s_E358_C1_H				  :std_logic_vector(11 downto 0) := x"2CC"; 
		s_E359_C1_H				  :std_logic_vector(11 downto 0) := x"2CE"; 
		s_E360_C1_H				  :std_logic_vector(11 downto 0) := x"2D0"; 
		s_E361_C1_H				  :std_logic_vector(11 downto 0) := x"2D2"; 
		s_E362_C1_H				  :std_logic_vector(11 downto 0) := x"2D4"; 
		s_E363_C1_H				  :std_logic_vector(11 downto 0) := x"2D6"; 
		s_E364_C1_H				  :std_logic_vector(11 downto 0) := x"2D8"; 
		s_E365_C1_H				  :std_logic_vector(11 downto 0) := x"2DA"; 
		s_E366_C1_H				  :std_logic_vector(11 downto 0) := x"2DC"; 
		s_E367_C1_H				  :std_logic_vector(11 downto 0) := x"2DE"; 
		s_E368_C1_H				  :std_logic_vector(11 downto 0) := x"2E0"; 
		s_E369_C1_H				  :std_logic_vector(11 downto 0) := x"2E2"; 
		s_E370_C1_H				  :std_logic_vector(11 downto 0) := x"2E4"; 
		s_E371_C1_H				  :std_logic_vector(11 downto 0) := x"2E6"; 
		s_E372_C1_H				  :std_logic_vector(11 downto 0) := x"2E8"; 
		s_E373_C1_H				  :std_logic_vector(11 downto 0) := x"2EA"; 
		s_E374_C1_H				  :std_logic_vector(11 downto 0) := x"2EC"; 
		s_E375_C1_H				  :std_logic_vector(11 downto 0) := x"2EE"; 
		s_E376_C1_H				  :std_logic_vector(11 downto 0) := x"2F0"; 
		s_E377_C1_H				  :std_logic_vector(11 downto 0) := x"2F2"; 
		s_E378_C1_H				  :std_logic_vector(11 downto 0) := x"2F4"; 
		s_E379_C1_H				  :std_logic_vector(11 downto 0) := x"2F6"; 
		s_E380_C1_H				  :std_logic_vector(11 downto 0) := x"2F8"; 
		s_E381_C1_H				  :std_logic_vector(11 downto 0) := x"2FA"; 
		s_E382_C1_H				  :std_logic_vector(11 downto 0) := x"2FC"; 
		s_E383_C1_H				  :std_logic_vector(11 downto 0) := x"2FE"; 
		s_E384_C1_H				  :std_logic_vector(11 downto 0) := x"300"; 
		s_E385_C1_H				  :std_logic_vector(11 downto 0) := x"302"; 
		s_E386_C1_H				  :std_logic_vector(11 downto 0) := x"304"; 
		s_E387_C1_H				  :std_logic_vector(11 downto 0) := x"306"; 
		s_E388_C1_H				  :std_logic_vector(11 downto 0) := x"308"; 
		s_E389_C1_H				  :std_logic_vector(11 downto 0) := x"30A"; 
		s_E390_C1_H				  :std_logic_vector(11 downto 0) := x"30C"; 
		s_E391_C1_H				  :std_logic_vector(11 downto 0) := x"30E"; 
		s_E392_C1_H				  :std_logic_vector(11 downto 0) := x"310"; 
		s_E393_C1_H				  :std_logic_vector(11 downto 0) := x"312"; 
		s_E394_C1_H				  :std_logic_vector(11 downto 0) := x"314"; 
		s_E395_C1_H				  :std_logic_vector(11 downto 0) := x"316"; 
		s_E396_C1_H				  :std_logic_vector(11 downto 0) := x"318"; 
		s_E397_C1_H				  :std_logic_vector(11 downto 0) := x"31A"; 
		s_E398_C1_H				  :std_logic_vector(11 downto 0) := x"31C"; 
		s_E399_C1_H				  :std_logic_vector(11 downto 0) := x"31E"; 
		s_E400_C1_H				  :std_logic_vector(11 downto 0) := x"320"; 
		s_E401_C1_H				  :std_logic_vector(11 downto 0) := x"322"; 
		s_E402_C1_H				  :std_logic_vector(11 downto 0) := x"324"; 
		s_E403_C1_H				  :std_logic_vector(11 downto 0) := x"326"; 
		s_E404_C1_H				  :std_logic_vector(11 downto 0) := x"328"; 
		s_E405_C1_H				  :std_logic_vector(11 downto 0) := x"32A"; 
		s_E406_C1_H				  :std_logic_vector(11 downto 0) := x"32C"; 
		s_E407_C1_H				  :std_logic_vector(11 downto 0) := x"32E"; 
		s_E408_C1_H				  :std_logic_vector(11 downto 0) := x"330"; 
		s_E409_C1_H				  :std_logic_vector(11 downto 0) := x"332"; 
		s_E410_C1_H				  :std_logic_vector(11 downto 0) := x"334"; 
		s_E411_C1_H				  :std_logic_vector(11 downto 0) := x"336"; 
		s_E412_C1_H				  :std_logic_vector(11 downto 0) := x"338"; 
		s_E413_C1_H				  :std_logic_vector(11 downto 0) := x"33A"; 
		s_E414_C1_H				  :std_logic_vector(11 downto 0) := x"33C"; 
		s_E415_C1_H				  :std_logic_vector(11 downto 0) := x"33E"; 
		s_E416_C1_H				  :std_logic_vector(11 downto 0) := x"340"; 
		s_E417_C1_H				  :std_logic_vector(11 downto 0) := x"342"; 
		s_E418_C1_H				  :std_logic_vector(11 downto 0) := x"344"; 
		s_E419_C1_H				  :std_logic_vector(11 downto 0) := x"346"; 
		s_E420_C1_H				  :std_logic_vector(11 downto 0) := x"348"; 
		s_E421_C1_H				  :std_logic_vector(11 downto 0) := x"34A"; 
		s_E422_C1_H				  :std_logic_vector(11 downto 0) := x"34C"; 
		s_E423_C1_H				  :std_logic_vector(11 downto 0) := x"34E"; 
		s_E424_C1_H				  :std_logic_vector(11 downto 0) := x"350"; 
		s_E425_C1_H				  :std_logic_vector(11 downto 0) := x"352"; 
		s_E426_C1_H				  :std_logic_vector(11 downto 0) := x"354"; 
		s_E427_C1_H				  :std_logic_vector(11 downto 0) := x"356"; 
		s_E428_C1_H				  :std_logic_vector(11 downto 0) := x"358"; 
		s_E429_C1_H				  :std_logic_vector(11 downto 0) := x"35A"; 
		s_E430_C1_H				  :std_logic_vector(11 downto 0) := x"35C"; 
		s_E431_C1_H				  :std_logic_vector(11 downto 0) := x"35E"; 
		s_E432_C1_H				  :std_logic_vector(11 downto 0) := x"360"; 
		s_E433_C1_H				  :std_logic_vector(11 downto 0) := x"362"; 
		s_E434_C1_H				  :std_logic_vector(11 downto 0) := x"364"; 
		s_E435_C1_H				  :std_logic_vector(11 downto 0) := x"366"; 
		s_E436_C1_H				  :std_logic_vector(11 downto 0) := x"368"; 
		s_E437_C1_H				  :std_logic_vector(11 downto 0) := x"36A"; 
		s_E438_C1_H				  :std_logic_vector(11 downto 0) := x"36C"; 
		s_E439_C1_H				  :std_logic_vector(11 downto 0) := x"36E"; 
		s_E440_C1_H				  :std_logic_vector(11 downto 0) := x"370"; 
		s_E441_C1_H				  :std_logic_vector(11 downto 0) := x"372"; 
		s_E442_C1_H				  :std_logic_vector(11 downto 0) := x"374"; 
		s_E443_C1_H				  :std_logic_vector(11 downto 0) := x"376"; 
		s_E444_C1_H				  :std_logic_vector(11 downto 0) := x"378"; 
		s_E445_C1_H				  :std_logic_vector(11 downto 0) := x"37A"; 
		s_E446_C1_H				  :std_logic_vector(11 downto 0) := x"37C"; 
		s_E447_C1_H				  :std_logic_vector(11 downto 0) := x"37E"; 
		s_E448_C1_H				  :std_logic_vector(11 downto 0) := x"380"; 
		s_E449_C1_H				  :std_logic_vector(11 downto 0) := x"382"; 
		s_E450_C1_H				  :std_logic_vector(11 downto 0) := x"384"; 
		s_E451_C1_H				  :std_logic_vector(11 downto 0) := x"386"; 
		s_E452_C1_H				  :std_logic_vector(11 downto 0) := x"388"; 
		s_E453_C1_H				  :std_logic_vector(11 downto 0) := x"38A"; 
		s_E454_C1_H				  :std_logic_vector(11 downto 0) := x"38C"; 
		s_E455_C1_H				  :std_logic_vector(11 downto 0) := x"38E"; 
		s_E456_C1_H				  :std_logic_vector(11 downto 0) := x"390"; 
		s_E457_C1_H				  :std_logic_vector(11 downto 0) := x"392"; 
		s_E458_C1_H				  :std_logic_vector(11 downto 0) := x"394"; 
		s_E459_C1_H				  :std_logic_vector(11 downto 0) := x"396"; 
		s_E460_C1_H				  :std_logic_vector(11 downto 0) := x"398"; 
		s_E461_C1_H				  :std_logic_vector(11 downto 0) := x"39A"; 
		s_E462_C1_H				  :std_logic_vector(11 downto 0) := x"39C"; 
		s_E463_C1_H				  :std_logic_vector(11 downto 0) := x"39E"; 
		s_E464_C1_H				  :std_logic_vector(11 downto 0) := x"3A0"; 
		s_E465_C1_H				  :std_logic_vector(11 downto 0) := x"3A2"; 
		s_E466_C1_H				  :std_logic_vector(11 downto 0) := x"3A4"; 
		s_E467_C1_H				  :std_logic_vector(11 downto 0) := x"3A6"; 
		s_E468_C1_H				  :std_logic_vector(11 downto 0) := x"3A8"; 
		s_E469_C1_H				  :std_logic_vector(11 downto 0) := x"3AA"; 
		s_E470_C1_H				  :std_logic_vector(11 downto 0) := x"3AC"; 
		s_E471_C1_H				  :std_logic_vector(11 downto 0) := x"3AE"; 
		s_E472_C1_H				  :std_logic_vector(11 downto 0) := x"3B0"; 
		s_E473_C1_H				  :std_logic_vector(11 downto 0) := x"3B2"; 
		s_E474_C1_H				  :std_logic_vector(11 downto 0) := x"3B4"; 
		s_E475_C1_H				  :std_logic_vector(11 downto 0) := x"3B6"; 
		s_E476_C1_H				  :std_logic_vector(11 downto 0) := x"3B8"; 
		s_E477_C1_H				  :std_logic_vector(11 downto 0) := x"3BA"; 
		s_E478_C1_H				  :std_logic_vector(11 downto 0) := x"3BC"; 
		s_E479_C1_H				  :std_logic_vector(11 downto 0) := x"3BE"; 
		s_E480_C1_H				  :std_logic_vector(11 downto 0) := x"3C0"; 
		s_E481_C1_H				  :std_logic_vector(11 downto 0) := x"3C2"; 
		s_E482_C1_H				  :std_logic_vector(11 downto 0) := x"3C4"; 
		s_E483_C1_H				  :std_logic_vector(11 downto 0) := x"3C6"; 
		s_E484_C1_H				  :std_logic_vector(11 downto 0) := x"3C8"; 
		s_E485_C1_H				  :std_logic_vector(11 downto 0) := x"3CA"; 
		s_E486_C1_H				  :std_logic_vector(11 downto 0) := x"3CC"; 
		s_E487_C1_H				  :std_logic_vector(11 downto 0) := x"3CE"; 
		s_E488_C1_H				  :std_logic_vector(11 downto 0) := x"3D0"; 
		s_E489_C1_H				  :std_logic_vector(11 downto 0) := x"3D2"; 
		s_E490_C1_H				  :std_logic_vector(11 downto 0) := x"3D4"; 
		s_E491_C1_H				  :std_logic_vector(11 downto 0) := x"3D6"; 
		s_E492_C1_H				  :std_logic_vector(11 downto 0) := x"3D8"; 
		s_E493_C1_H				  :std_logic_vector(11 downto 0) := x"3DA"; 
		s_E494_C1_H				  :std_logic_vector(11 downto 0) := x"3DC"; 
		s_E495_C1_H				  :std_logic_vector(11 downto 0) := x"3DE"; 
		s_E496_C1_H				  :std_logic_vector(11 downto 0) := x"3E0"; 
		s_E497_C1_H				  :std_logic_vector(11 downto 0) := x"3E2"; 
		s_E498_C1_H				  :std_logic_vector(11 downto 0) := x"3E4"; 
		s_E499_C1_H				  :std_logic_vector(11 downto 0) := x"3E6"; 
		s_E500_C1_H				  :std_logic_vector(11 downto 0) := x"3E8"; 
		s_E501_C1_H				  :std_logic_vector(11 downto 0) := x"3EA"; 
		s_E502_C1_H				  :std_logic_vector(11 downto 0) := x"3EC"; 
		s_E503_C1_H				  :std_logic_vector(11 downto 0) := x"3EE"; 
		s_E504_C1_H				  :std_logic_vector(11 downto 0) := x"3F0"; 
		s_E505_C1_H				  :std_logic_vector(11 downto 0) := x"3F2"; 
		s_E506_C1_H				  :std_logic_vector(11 downto 0) := x"3F4"; 
		s_E507_C1_H				  :std_logic_vector(11 downto 0) := x"3F6"; 
		s_E508_C1_H				  :std_logic_vector(11 downto 0) := x"3F8"; 
		s_E509_C1_H				  :std_logic_vector(11 downto 0) := x"3FA"; 
		s_E510_C1_H				  :std_logic_vector(11 downto 0) := x"3FC"; 
		s_E511_C1_H				  :std_logic_vector(11 downto 0) := x"3FE"; 
		s_E512_C1_H				  :std_logic_vector(11 downto 0) := x"400"; 
		s_E513_C1_H				  :std_logic_vector(11 downto 0) := x"402"; 
		s_E514_C1_H				  :std_logic_vector(11 downto 0) := x"404"; 
		s_E515_C1_H				  :std_logic_vector(11 downto 0) := x"406"; 
		s_E516_C1_H				  :std_logic_vector(11 downto 0) := x"408"; 
		s_E517_C1_H				  :std_logic_vector(11 downto 0) := x"40A"; 
		s_E518_C1_H				  :std_logic_vector(11 downto 0) := x"40C"; 
		s_E519_C1_H				  :std_logic_vector(11 downto 0) := x"40E"; 
		s_E520_C1_H				  :std_logic_vector(11 downto 0) := x"410"; 
		s_E521_C1_H				  :std_logic_vector(11 downto 0) := x"412"; 
		s_E522_C1_H				  :std_logic_vector(11 downto 0) := x"414"; 
		s_E523_C1_H				  :std_logic_vector(11 downto 0) := x"416"; 
		s_E524_C1_H				  :std_logic_vector(11 downto 0) := x"418"; 
		s_E525_C1_H				  :std_logic_vector(11 downto 0) := x"41A"; 
		s_E526_C1_H				  :std_logic_vector(11 downto 0) := x"41C"; 
		s_E527_C1_H				  :std_logic_vector(11 downto 0) := x"41E"; 
		s_E528_C1_H				  :std_logic_vector(11 downto 0) := x"420"; 
		s_E529_C1_H				  :std_logic_vector(11 downto 0) := x"422"; 
		s_E530_C1_H				  :std_logic_vector(11 downto 0) := x"424"; 
		s_E531_C1_H				  :std_logic_vector(11 downto 0) := x"426"; 
		s_E532_C1_H				  :std_logic_vector(11 downto 0) := x"428"; 
		s_E533_C1_H				  :std_logic_vector(11 downto 0) := x"42A"; 
		s_E534_C1_H				  :std_logic_vector(11 downto 0) := x"42C"; 
		s_E535_C1_H				  :std_logic_vector(11 downto 0) := x"42E"; 
		s_E536_C1_H				  :std_logic_vector(11 downto 0) := x"430"; 
		s_E537_C1_H				  :std_logic_vector(11 downto 0) := x"432"; 
		s_E538_C1_H				  :std_logic_vector(11 downto 0) := x"434"; 
		s_E539_C1_H				  :std_logic_vector(11 downto 0) := x"436"; 
		s_E540_C1_H				  :std_logic_vector(11 downto 0) := x"438"; 
		s_E541_C1_H				  :std_logic_vector(11 downto 0) := x"43A"; 
		s_E542_C1_H				  :std_logic_vector(11 downto 0) := x"43C"; 
		s_E543_C1_H				  :std_logic_vector(11 downto 0) := x"43E"; 
		s_E544_C1_H				  :std_logic_vector(11 downto 0) := x"440"; 
		s_E545_C1_H				  :std_logic_vector(11 downto 0) := x"442"; 
		s_E546_C1_H				  :std_logic_vector(11 downto 0) := x"444"; 
		s_E547_C1_H				  :std_logic_vector(11 downto 0) := x"446"; 
		s_E548_C1_H				  :std_logic_vector(11 downto 0) := x"448"; 
		s_E549_C1_H				  :std_logic_vector(11 downto 0) := x"44A"; 
		s_E550_C1_H				  :std_logic_vector(11 downto 0) := x"44C"; 
		s_E551_C1_H				  :std_logic_vector(11 downto 0) := x"44E"; 
		s_E552_C1_H				  :std_logic_vector(11 downto 0) := x"450"; 
		s_E553_C1_H				  :std_logic_vector(11 downto 0) := x"452"; 
		s_E554_C1_H				  :std_logic_vector(11 downto 0) := x"454"; 
		s_E555_C1_H				  :std_logic_vector(11 downto 0) := x"456"; 
		s_E556_C1_H				  :std_logic_vector(11 downto 0) := x"458"; 
		s_E557_C1_H				  :std_logic_vector(11 downto 0) := x"45A"; 
		s_E558_C1_H				  :std_logic_vector(11 downto 0) := x"45C"; 
		s_E559_C1_H				  :std_logic_vector(11 downto 0) := x"45E"; 
		s_E560_C1_H				  :std_logic_vector(11 downto 0) := x"460"; 
		s_E561_C1_H				  :std_logic_vector(11 downto 0) := x"462"; 
		s_E562_C1_H				  :std_logic_vector(11 downto 0) := x"464"; 
		s_E563_C1_H				  :std_logic_vector(11 downto 0) := x"466"; 
		s_E564_C1_H				  :std_logic_vector(11 downto 0) := x"468"; 
		s_E565_C1_H				  :std_logic_vector(11 downto 0) := x"46A"; 
		s_E566_C1_H				  :std_logic_vector(11 downto 0) := x"46C"; 
		s_E567_C1_H				  :std_logic_vector(11 downto 0) := x"46E"; 
		s_E568_C1_H				  :std_logic_vector(11 downto 0) := x"470"; 
		s_E569_C1_H				  :std_logic_vector(11 downto 0) := x"472"; 
		s_E570_C1_H				  :std_logic_vector(11 downto 0) := x"474"; 
		s_E571_C1_H				  :std_logic_vector(11 downto 0) := x"476"; 
		s_E572_C1_H				  :std_logic_vector(11 downto 0) := x"478"; 
		s_E573_C1_H				  :std_logic_vector(11 downto 0) := x"47A"; 
		s_E574_C1_H				  :std_logic_vector(11 downto 0) := x"47C"; 
		s_E575_C1_H				  :std_logic_vector(11 downto 0) := x"47E"; 
		s_E576_C1_H				  :std_logic_vector(11 downto 0) := x"480"; 
		s_E577_C1_H				  :std_logic_vector(11 downto 0) := x"482"; 
		s_E578_C1_H				  :std_logic_vector(11 downto 0) := x"484"; 
		s_E579_C1_H				  :std_logic_vector(11 downto 0) := x"486"; 
		s_E580_C1_H				  :std_logic_vector(11 downto 0) := x"488"; 
		s_E581_C1_H				  :std_logic_vector(11 downto 0) := x"48A"; 
		s_E582_C1_H				  :std_logic_vector(11 downto 0) := x"48C"; 
		s_E583_C1_H				  :std_logic_vector(11 downto 0) := x"48E"; 
		s_E584_C1_H				  :std_logic_vector(11 downto 0) := x"490"; 
		s_E585_C1_H				  :std_logic_vector(11 downto 0) := x"492"; 
		s_E586_C1_H				  :std_logic_vector(11 downto 0) := x"494"; 
		s_E587_C1_H				  :std_logic_vector(11 downto 0) := x"496"; 
		s_E588_C1_H				  :std_logic_vector(11 downto 0) := x"498"; 
		s_E589_C1_H				  :std_logic_vector(11 downto 0) := x"49A"; 
		s_E590_C1_H				  :std_logic_vector(11 downto 0) := x"49C"; 
		s_E591_C1_H				  :std_logic_vector(11 downto 0) := x"49E"; 
		s_E592_C1_H				  :std_logic_vector(11 downto 0) := x"4A0"; 
		s_E593_C1_H				  :std_logic_vector(11 downto 0) := x"4A2"; 
		s_E594_C1_H				  :std_logic_vector(11 downto 0) := x"4A4"; 
		s_E595_C1_H				  :std_logic_vector(11 downto 0) := x"4A6"; 
		s_E596_C1_H				  :std_logic_vector(11 downto 0) := x"4A8"; 
		s_E597_C1_H				  :std_logic_vector(11 downto 0) := x"4AA"; 
		s_E598_C1_H				  :std_logic_vector(11 downto 0) := x"4AC"; 
		s_E599_C1_H				  :std_logic_vector(11 downto 0) := x"4AE"; 
		s_E600_C1_H				  :std_logic_vector(11 downto 0) := x"4B0"; 
		s_E601_C1_H				  :std_logic_vector(11 downto 0) := x"4B2"; 
		s_E602_C1_H				  :std_logic_vector(11 downto 0) := x"4B4"; 
		s_E603_C1_H				  :std_logic_vector(11 downto 0) := x"4B6"; 
		s_E604_C1_H				  :std_logic_vector(11 downto 0) := x"4B8"; 
		s_E605_C1_H				  :std_logic_vector(11 downto 0) := x"4BA"; 
		s_E606_C1_H				  :std_logic_vector(11 downto 0) := x"4BC"; 
		s_E607_C1_H				  :std_logic_vector(11 downto 0) := x"4BE"; 
		s_E608_C1_H				  :std_logic_vector(11 downto 0) := x"4C0"; 
		s_E609_C1_H				  :std_logic_vector(11 downto 0) := x"4C2"; 
		s_E610_C1_H				  :std_logic_vector(11 downto 0) := x"4C4"; 
		s_E611_C1_H				  :std_logic_vector(11 downto 0) := x"4C6"; 
		s_E612_C1_H				  :std_logic_vector(11 downto 0) := x"4C8"; 
		s_E613_C1_H				  :std_logic_vector(11 downto 0) := x"4CA"; 
		s_E614_C1_H				  :std_logic_vector(11 downto 0) := x"4CC"; 
		s_E615_C1_H				  :std_logic_vector(11 downto 0) := x"4CE"; 
		s_E616_C1_H				  :std_logic_vector(11 downto 0) := x"4D0"; 
		s_E617_C1_H				  :std_logic_vector(11 downto 0) := x"4D2"; 
		s_E618_C1_H				  :std_logic_vector(11 downto 0) := x"4D4"; 
		s_E619_C1_H				  :std_logic_vector(11 downto 0) := x"4D6"; 
		s_E620_C1_H				  :std_logic_vector(11 downto 0) := x"4D8"; 
		s_E621_C1_H				  :std_logic_vector(11 downto 0) := x"4DA"; 
		s_E622_C1_H				  :std_logic_vector(11 downto 0) := x"4DC"; 
		s_E623_C1_H				  :std_logic_vector(11 downto 0) := x"4DE"; 
		s_E624_C1_H				  :std_logic_vector(11 downto 0) := x"4E0"; 
		s_E625_C1_H				  :std_logic_vector(11 downto 0) := x"4E2"; 
		s_E626_C1_H				  :std_logic_vector(11 downto 0) := x"4E4"; 
		s_E627_C1_H				  :std_logic_vector(11 downto 0) := x"4E6"; 
		s_E628_C1_H				  :std_logic_vector(11 downto 0) := x"4E8"; 
		s_E629_C1_H				  :std_logic_vector(11 downto 0) := x"4EA"; 
		s_E630_C1_H				  :std_logic_vector(11 downto 0) := x"4EC"; 
		s_E631_C1_H				  :std_logic_vector(11 downto 0) := x"4EE"; 
		s_E632_C1_H				  :std_logic_vector(11 downto 0) := x"4F0"; 
		s_E633_C1_H				  :std_logic_vector(11 downto 0) := x"4F2"; 
		s_E634_C1_H				  :std_logic_vector(11 downto 0) := x"4F4"; 
		s_E635_C1_H				  :std_logic_vector(11 downto 0) := x"4F6"; 
		s_E636_C1_H				  :std_logic_vector(11 downto 0) := x"4F8"; 
		s_E637_C1_H				  :std_logic_vector(11 downto 0) := x"4FA"; 
		s_E638_C1_H				  :std_logic_vector(11 downto 0) := x"4FC"; 
		s_E639_C1_H				  :std_logic_vector(11 downto 0) := x"4FE"; 
		s_E640_C1_H				  :std_logic_vector(11 downto 0) := x"500"; 
		s_E641_C1_H				  :std_logic_vector(11 downto 0) := x"502"; 
		s_E642_C1_H				  :std_logic_vector(11 downto 0) := x"504"; 
		s_E643_C1_H				  :std_logic_vector(11 downto 0) := x"506"; 
		s_E644_C1_H				  :std_logic_vector(11 downto 0) := x"508"; 
		s_E645_C1_H				  :std_logic_vector(11 downto 0) := x"50A"; 
		s_E646_C1_H				  :std_logic_vector(11 downto 0) := x"50C"; 
		s_E647_C1_H				  :std_logic_vector(11 downto 0) := x"50E"; 
		s_E648_C1_H				  :std_logic_vector(11 downto 0) := x"510"; 
		s_E649_C1_H				  :std_logic_vector(11 downto 0) := x"512"; 
		s_E650_C1_H				  :std_logic_vector(11 downto 0) := x"514"; 
		s_E651_C1_H				  :std_logic_vector(11 downto 0) := x"516"; 
		s_E652_C1_H				  :std_logic_vector(11 downto 0) := x"518"; 
		s_E653_C1_H				  :std_logic_vector(11 downto 0) := x"51A"; 
		s_E654_C1_H				  :std_logic_vector(11 downto 0) := x"51C"; 
		s_E655_C1_H				  :std_logic_vector(11 downto 0) := x"51E"; 
		s_E656_C1_H				  :std_logic_vector(11 downto 0) := x"520"; 
		s_E657_C1_H				  :std_logic_vector(11 downto 0) := x"522"; 
		s_E658_C1_H				  :std_logic_vector(11 downto 0) := x"524"; 
		s_E659_C1_H				  :std_logic_vector(11 downto 0) := x"526"; 
		s_E660_C1_H				  :std_logic_vector(11 downto 0) := x"528"; 
		s_E661_C1_H				  :std_logic_vector(11 downto 0) := x"52A"; 
		s_E662_C1_H				  :std_logic_vector(11 downto 0) := x"52C"; 
		s_E663_C1_H				  :std_logic_vector(11 downto 0) := x"52E"; 
		s_E664_C1_H				  :std_logic_vector(11 downto 0) := x"530"; 
		s_E665_C1_H				  :std_logic_vector(11 downto 0) := x"532"; 
		s_E666_C1_H				  :std_logic_vector(11 downto 0) := x"534"; 
		s_E667_C1_H				  :std_logic_vector(11 downto 0) := x"536"; 
		s_E668_C1_H				  :std_logic_vector(11 downto 0) := x"538"; 
		s_E669_C1_H				  :std_logic_vector(11 downto 0) := x"53A"; 
		s_E670_C1_H				  :std_logic_vector(11 downto 0) := x"53C"; 
		s_E671_C1_H				  :std_logic_vector(11 downto 0) := x"53E"; 
		s_E672_C1_H				  :std_logic_vector(11 downto 0) := x"540"; 
		s_E673_C1_H				  :std_logic_vector(11 downto 0) := x"542"; 
		s_E674_C1_H				  :std_logic_vector(11 downto 0) := x"544"; 
		s_E675_C1_H				  :std_logic_vector(11 downto 0) := x"546"; 
		s_E676_C1_H				  :std_logic_vector(11 downto 0) := x"548"; 
		s_E677_C1_H				  :std_logic_vector(11 downto 0) := x"54A"; 
		s_E678_C1_H				  :std_logic_vector(11 downto 0) := x"54C"; 
		s_E679_C1_H				  :std_logic_vector(11 downto 0) := x"54E"; 
		s_E680_C1_H				  :std_logic_vector(11 downto 0) := x"550"; 
		s_E681_C1_H				  :std_logic_vector(11 downto 0) := x"552"; 
		s_E682_C1_H				  :std_logic_vector(11 downto 0) := x"554"; 
		s_E683_C1_H				  :std_logic_vector(11 downto 0) := x"556"; 
		s_E684_C1_H				  :std_logic_vector(11 downto 0) := x"558"; 
		s_E685_C1_H				  :std_logic_vector(11 downto 0) := x"55A"; 
		s_E686_C1_H				  :std_logic_vector(11 downto 0) := x"55C"; 
		s_E687_C1_H				  :std_logic_vector(11 downto 0) := x"55E"; 
		s_E688_C1_H				  :std_logic_vector(11 downto 0) := x"560"; 
		s_E689_C1_H				  :std_logic_vector(11 downto 0) := x"562"; 
		s_E690_C1_H				  :std_logic_vector(11 downto 0) := x"564"; 
		s_E691_C1_H				  :std_logic_vector(11 downto 0) := x"566"; 
		s_E692_C1_H				  :std_logic_vector(11 downto 0) := x"568"; 
		s_E693_C1_H				  :std_logic_vector(11 downto 0) := x"56A"; 
		s_E694_C1_H				  :std_logic_vector(11 downto 0) := x"56C"; 
		s_E695_C1_H				  :std_logic_vector(11 downto 0) := x"56E"; 
		s_E696_C1_H				  :std_logic_vector(11 downto 0) := x"570"; 
		s_E697_C1_H				  :std_logic_vector(11 downto 0) := x"572"; 
		s_E698_C1_H				  :std_logic_vector(11 downto 0) := x"574"; 
		s_E699_C1_H				  :std_logic_vector(11 downto 0) := x"576"; 
		s_E700_C1_H				  :std_logic_vector(11 downto 0) := x"578"; 
		s_E701_C1_H				  :std_logic_vector(11 downto 0) := x"57A"; 
		s_E702_C1_H				  :std_logic_vector(11 downto 0) := x"57C"; 
		s_E703_C1_H				  :std_logic_vector(11 downto 0) := x"57E"; 
		s_E704_C1_H				  :std_logic_vector(11 downto 0) := x"580"; 
		s_E705_C1_H				  :std_logic_vector(11 downto 0) := x"582"; 
		s_E706_C1_H				  :std_logic_vector(11 downto 0) := x"584"; 
		s_E707_C1_H				  :std_logic_vector(11 downto 0) := x"586"; 
		s_E708_C1_H				  :std_logic_vector(11 downto 0) := x"588"; 
		s_E709_C1_H				  :std_logic_vector(11 downto 0) := x"58A"; 
		s_E710_C1_H				  :std_logic_vector(11 downto 0) := x"58C"; 
		s_E711_C1_H				  :std_logic_vector(11 downto 0) := x"58E"; 
		s_E712_C1_H				  :std_logic_vector(11 downto 0) := x"590"; 
		s_E713_C1_H				  :std_logic_vector(11 downto 0) := x"592"; 
		s_E714_C1_H				  :std_logic_vector(11 downto 0) := x"594"; 
		s_E715_C1_H				  :std_logic_vector(11 downto 0) := x"596"; 
		s_E716_C1_H				  :std_logic_vector(11 downto 0) := x"598"; 
		s_E717_C1_H				  :std_logic_vector(11 downto 0) := x"59A"; 
		s_E718_C1_H				  :std_logic_vector(11 downto 0) := x"59C"; 
		s_E719_C1_H				  :std_logic_vector(11 downto 0) := x"59E"; 
		s_E720_C1_H				  :std_logic_vector(11 downto 0) := x"5A0"; 
		s_E721_C1_H				  :std_logic_vector(11 downto 0) := x"5A2"; 
		s_E722_C1_H				  :std_logic_vector(11 downto 0) := x"5A4"; 
		s_E723_C1_H				  :std_logic_vector(11 downto 0) := x"5A6"; 
		s_E724_C1_H				  :std_logic_vector(11 downto 0) := x"5A8"; 
		s_E725_C1_H				  :std_logic_vector(11 downto 0) := x"5AA"; 
		s_E726_C1_H				  :std_logic_vector(11 downto 0) := x"5AC"; 
		s_E727_C1_H				  :std_logic_vector(11 downto 0) := x"5AE"; 
		s_E728_C1_H				  :std_logic_vector(11 downto 0) := x"5B0"; 
		s_E729_C1_H				  :std_logic_vector(11 downto 0) := x"5B2"; 
		s_E730_C1_H				  :std_logic_vector(11 downto 0) := x"5B4"; 
		s_E731_C1_H				  :std_logic_vector(11 downto 0) := x"5B6"; 
		s_E732_C1_H				  :std_logic_vector(11 downto 0) := x"5B8"; 
		s_E733_C1_H				  :std_logic_vector(11 downto 0) := x"5BA"; 
		s_E734_C1_H				  :std_logic_vector(11 downto 0) := x"5BC"; 
		s_E735_C1_H				  :std_logic_vector(11 downto 0) := x"5BE"; 
		s_E736_C1_H				  :std_logic_vector(11 downto 0) := x"5C0"; 
		s_E737_C1_H				  :std_logic_vector(11 downto 0) := x"5C2"; 
		s_E738_C1_H				  :std_logic_vector(11 downto 0) := x"5C4"; 
		s_E739_C1_H				  :std_logic_vector(11 downto 0) := x"5C6"; 
		s_E740_C1_H				  :std_logic_vector(11 downto 0) := x"5C8"; 
		s_E741_C1_H				  :std_logic_vector(11 downto 0) := x"5CA"; 
		s_E742_C1_H				  :std_logic_vector(11 downto 0) := x"5CC"; 
		s_E743_C1_H				  :std_logic_vector(11 downto 0) := x"5CE"; 
		s_E744_C1_H				  :std_logic_vector(11 downto 0) := x"5D0"; 
		s_E745_C1_H				  :std_logic_vector(11 downto 0) := x"5D2"; 
		s_E746_C1_H				  :std_logic_vector(11 downto 0) := x"5D4"; 
		s_E747_C1_H				  :std_logic_vector(11 downto 0) := x"5D6"; 
		s_E748_C1_H				  :std_logic_vector(11 downto 0) := x"5D8"; 
		s_E749_C1_H				  :std_logic_vector(11 downto 0) := x"5DA"; 
		s_E750_C1_H				  :std_logic_vector(11 downto 0) := x"5DC"; 
		s_E751_C1_H				  :std_logic_vector(11 downto 0) := x"5DE"; 
		s_E752_C1_H				  :std_logic_vector(11 downto 0) := x"5E0"; 
		s_E753_C1_H				  :std_logic_vector(11 downto 0) := x"5E2"; 
		s_E754_C1_H				  :std_logic_vector(11 downto 0) := x"5E4"; 
		s_E755_C1_H				  :std_logic_vector(11 downto 0) := x"5E6"; 
		s_E756_C1_H				  :std_logic_vector(11 downto 0) := x"5E8"; 
		s_E757_C1_H				  :std_logic_vector(11 downto 0) := x"5EA"; 
		s_E758_C1_H				  :std_logic_vector(11 downto 0) := x"5EC"; 
		s_E759_C1_H				  :std_logic_vector(11 downto 0) := x"5EE"; 
		s_E760_C1_H				  :std_logic_vector(11 downto 0) := x"5F0"; 
		s_E761_C1_H				  :std_logic_vector(11 downto 0) := x"5F2"; 
		s_E762_C1_H				  :std_logic_vector(11 downto 0) := x"5F4"; 
		s_E763_C1_H				  :std_logic_vector(11 downto 0) := x"5F6"; 
		s_E764_C1_H				  :std_logic_vector(11 downto 0) := x"5F8"; 
		s_E765_C1_H				  :std_logic_vector(11 downto 0) := x"5FA"; 
		s_E766_C1_H				  :std_logic_vector(11 downto 0) := x"5FC"; 
		s_E767_C1_H				  :std_logic_vector(11 downto 0) := x"5FE"; 
		s_E768_C1_H				  :std_logic_vector(11 downto 0) := x"600"; 
		s_E769_C1_H				  :std_logic_vector(11 downto 0) := x"602"; 
		s_E770_C1_H				  :std_logic_vector(11 downto 0) := x"604"; 
		s_E771_C1_H				  :std_logic_vector(11 downto 0) := x"606"; 
		s_E772_C1_H				  :std_logic_vector(11 downto 0) := x"608"; 
		s_E773_C1_H				  :std_logic_vector(11 downto 0) := x"60A"; 
		s_E774_C1_H				  :std_logic_vector(11 downto 0) := x"60C"; 
		s_E775_C1_H				  :std_logic_vector(11 downto 0) := x"60E"; 
		s_E776_C1_H				  :std_logic_vector(11 downto 0) := x"610"; 
		s_E777_C1_H				  :std_logic_vector(11 downto 0) := x"612"; 
		s_E778_C1_H				  :std_logic_vector(11 downto 0) := x"614"; 
		s_E779_C1_H				  :std_logic_vector(11 downto 0) := x"616"; 
		s_E780_C1_H				  :std_logic_vector(11 downto 0) := x"618"; 
		s_E781_C1_H				  :std_logic_vector(11 downto 0) := x"61A"; 
		s_E782_C1_H				  :std_logic_vector(11 downto 0) := x"61C"; 
		s_E783_C1_H				  :std_logic_vector(11 downto 0) := x"61E"; 
		s_E784_C1_H				  :std_logic_vector(11 downto 0) := x"620"; 
		s_E785_C1_H				  :std_logic_vector(11 downto 0) := x"622"; 
		s_E786_C1_H				  :std_logic_vector(11 downto 0) := x"624"; 
		s_E787_C1_H				  :std_logic_vector(11 downto 0) := x"626"; 
		s_E788_C1_H				  :std_logic_vector(11 downto 0) := x"628"; 
		s_E789_C1_H				  :std_logic_vector(11 downto 0) := x"62A"; 
		s_E790_C1_H				  :std_logic_vector(11 downto 0) := x"62C"; 
		s_E791_C1_H				  :std_logic_vector(11 downto 0) := x"62E"; 
		s_E792_C1_H				  :std_logic_vector(11 downto 0) := x"630"; 
		s_E793_C1_H				  :std_logic_vector(11 downto 0) := x"632"; 
		s_E794_C1_H				  :std_logic_vector(11 downto 0) := x"634"; 
		s_E795_C1_H				  :std_logic_vector(11 downto 0) := x"636"; 
		s_E796_C1_H				  :std_logic_vector(11 downto 0) := x"638"; 
		s_E797_C1_H				  :std_logic_vector(11 downto 0) := x"63A"; 
		s_E798_C1_H				  :std_logic_vector(11 downto 0) := x"63C"; 
		s_E799_C1_H				  :std_logic_vector(11 downto 0) := x"63E"; 
		s_E800_C1_H				  :std_logic_vector(11 downto 0) := x"640"; 
		s_E801_C1_H				  :std_logic_vector(11 downto 0) := x"642"; 
		s_E802_C1_H				  :std_logic_vector(11 downto 0) := x"644"; 
		s_E803_C1_H				  :std_logic_vector(11 downto 0) := x"646"; 
		s_E804_C1_H				  :std_logic_vector(11 downto 0) := x"648"; 
		s_E805_C1_H				  :std_logic_vector(11 downto 0) := x"64A"; 
		s_E806_C1_H				  :std_logic_vector(11 downto 0) := x"64C"; 
		s_E807_C1_H				  :std_logic_vector(11 downto 0) := x"64E"; 
		s_E808_C1_H				  :std_logic_vector(11 downto 0) := x"650"; 
		s_E809_C1_H				  :std_logic_vector(11 downto 0) := x"652"; 
		s_E810_C1_H				  :std_logic_vector(11 downto 0) := x"654"; 
		s_E811_C1_H				  :std_logic_vector(11 downto 0) := x"656"; 
		s_E812_C1_H				  :std_logic_vector(11 downto 0) := x"658"; 
		s_E813_C1_H				  :std_logic_vector(11 downto 0) := x"65A"; 
		s_E814_C1_H				  :std_logic_vector(11 downto 0) := x"65C"; 
		s_E815_C1_H				  :std_logic_vector(11 downto 0) := x"65E"; 
		s_E816_C1_H				  :std_logic_vector(11 downto 0) := x"660"; 
		s_E817_C1_H				  :std_logic_vector(11 downto 0) := x"662"; 
		s_E818_C1_H				  :std_logic_vector(11 downto 0) := x"664"; 
		s_E819_C1_H				  :std_logic_vector(11 downto 0) := x"666"; 
		s_E820_C1_H				  :std_logic_vector(11 downto 0) := x"668"; 
		s_E821_C1_H				  :std_logic_vector(11 downto 0) := x"66A"; 
		s_E822_C1_H				  :std_logic_vector(11 downto 0) := x"66C"; 
		s_E823_C1_H				  :std_logic_vector(11 downto 0) := x"66E"; 
		s_E824_C1_H				  :std_logic_vector(11 downto 0) := x"670"; 
		s_E825_C1_H				  :std_logic_vector(11 downto 0) := x"672"; 
		s_E826_C1_H				  :std_logic_vector(11 downto 0) := x"674"; 
		s_E827_C1_H				  :std_logic_vector(11 downto 0) := x"676"; 
		s_E828_C1_H				  :std_logic_vector(11 downto 0) := x"678"; 
		s_E829_C1_H				  :std_logic_vector(11 downto 0) := x"67A"; 
		s_E830_C1_H				  :std_logic_vector(11 downto 0) := x"67C"; 
		s_E831_C1_H				  :std_logic_vector(11 downto 0) := x"67E"; 
		s_E832_C1_H				  :std_logic_vector(11 downto 0) := x"680"; 
		s_E833_C1_H				  :std_logic_vector(11 downto 0) := x"682"; 
		s_E834_C1_H				  :std_logic_vector(11 downto 0) := x"684"; 
		s_E835_C1_H				  :std_logic_vector(11 downto 0) := x"686"; 
		s_E836_C1_H				  :std_logic_vector(11 downto 0) := x"688"; 
		s_E837_C1_H				  :std_logic_vector(11 downto 0) := x"68A"; 
		s_E838_C1_H				  :std_logic_vector(11 downto 0) := x"68C"; 
		s_E839_C1_H				  :std_logic_vector(11 downto 0) := x"68E"; 
		s_E840_C1_H				  :std_logic_vector(11 downto 0) := x"690"; 
		s_E841_C1_H				  :std_logic_vector(11 downto 0) := x"692"; 
		s_E842_C1_H				  :std_logic_vector(11 downto 0) := x"694"; 
		s_E843_C1_H				  :std_logic_vector(11 downto 0) := x"696"; 
		s_E844_C1_H				  :std_logic_vector(11 downto 0) := x"698"; 
		s_E845_C1_H				  :std_logic_vector(11 downto 0) := x"69A"; 
		s_E846_C1_H				  :std_logic_vector(11 downto 0) := x"69C"; 
		s_E847_C1_H				  :std_logic_vector(11 downto 0) := x"69E"; 
		s_E848_C1_H				  :std_logic_vector(11 downto 0) := x"6A0"; 
		s_E849_C1_H				  :std_logic_vector(11 downto 0) := x"6A2"; 
		s_E850_C1_H				  :std_logic_vector(11 downto 0) := x"6A4"; 
		s_E851_C1_H				  :std_logic_vector(11 downto 0) := x"6A6"; 
		s_E852_C1_H				  :std_logic_vector(11 downto 0) := x"6A8"; 
		s_E853_C1_H				  :std_logic_vector(11 downto 0) := x"6AA"; 
		s_E854_C1_H				  :std_logic_vector(11 downto 0) := x"6AC"; 
		s_E855_C1_H				  :std_logic_vector(11 downto 0) := x"6AE"; 
		s_E856_C1_H				  :std_logic_vector(11 downto 0) := x"6B0"; 
		s_E857_C1_H				  :std_logic_vector(11 downto 0) := x"6B2"; 
		s_E858_C1_H				  :std_logic_vector(11 downto 0) := x"6B4"; 
		s_E859_C1_H				  :std_logic_vector(11 downto 0) := x"6B6"; 
		s_E860_C1_H				  :std_logic_vector(11 downto 0) := x"6B8"; 
		s_E861_C1_H				  :std_logic_vector(11 downto 0) := x"6BA"; 
		s_E862_C1_H				  :std_logic_vector(11 downto 0) := x"6BC"; 
		s_E863_C1_H				  :std_logic_vector(11 downto 0) := x"6BE"; 
		s_E864_C1_H				  :std_logic_vector(11 downto 0) := x"6C0"; 
		s_E865_C1_H				  :std_logic_vector(11 downto 0) := x"6C2"; 
		s_E866_C1_H				  :std_logic_vector(11 downto 0) := x"6C4"; 
		s_E867_C1_H				  :std_logic_vector(11 downto 0) := x"6C6"; 
		s_E868_C1_H				  :std_logic_vector(11 downto 0) := x"6C8"; 
		s_E869_C1_H				  :std_logic_vector(11 downto 0) := x"6CA"; 
		s_E870_C1_H				  :std_logic_vector(11 downto 0) := x"6CC"; 
		s_E871_C1_H				  :std_logic_vector(11 downto 0) := x"6CE"; 
		s_E872_C1_H				  :std_logic_vector(11 downto 0) := x"6D0"; 
		s_E873_C1_H				  :std_logic_vector(11 downto 0) := x"6D2"; 
		s_E874_C1_H				  :std_logic_vector(11 downto 0) := x"6D4"; 
		s_E875_C1_H				  :std_logic_vector(11 downto 0) := x"6D6"; 
		s_E876_C1_H				  :std_logic_vector(11 downto 0) := x"6D8"; 
		s_E877_C1_H				  :std_logic_vector(11 downto 0) := x"6DA"; 
		s_E878_C1_H				  :std_logic_vector(11 downto 0) := x"6DC"; 
		s_E879_C1_H				  :std_logic_vector(11 downto 0) := x"6DE"; 
		s_E880_C1_H				  :std_logic_vector(11 downto 0) := x"6E0"; 
		s_E881_C1_H				  :std_logic_vector(11 downto 0) := x"6E2"; 
		s_E882_C1_H				  :std_logic_vector(11 downto 0) := x"6E4"; 
		s_E883_C1_H				  :std_logic_vector(11 downto 0) := x"6E6"; 
		s_E884_C1_H				  :std_logic_vector(11 downto 0) := x"6E8"; 
		s_E885_C1_H				  :std_logic_vector(11 downto 0) := x"6EA"; 
		s_E886_C1_H				  :std_logic_vector(11 downto 0) := x"6EC"; 
		s_E887_C1_H				  :std_logic_vector(11 downto 0) := x"6EE"; 
		s_E888_C1_H				  :std_logic_vector(11 downto 0) := x"6F0"; 
		s_E889_C1_H				  :std_logic_vector(11 downto 0) := x"6F2"; 
		s_E890_C1_H				  :std_logic_vector(11 downto 0) := x"6F4"; 
		s_E891_C1_H				  :std_logic_vector(11 downto 0) := x"6F6"; 
		s_E892_C1_H				  :std_logic_vector(11 downto 0) := x"6F8"; 
		s_E893_C1_H				  :std_logic_vector(11 downto 0) := x"6FA"; 
		s_E894_C1_H				  :std_logic_vector(11 downto 0) := x"6FC"; 
		s_E895_C1_H				  :std_logic_vector(11 downto 0) := x"6FE"; 
		s_E896_C1_H				  :std_logic_vector(11 downto 0) := x"700"; 
		s_E897_C1_H				  :std_logic_vector(11 downto 0) := x"702"; 
		s_E898_C1_H				  :std_logic_vector(11 downto 0) := x"704"; 
		s_E899_C1_H				  :std_logic_vector(11 downto 0) := x"706"; 
		s_E900_C1_H				  :std_logic_vector(11 downto 0) := x"708"; 
		s_E901_C1_H				  :std_logic_vector(11 downto 0) := x"70A"; 
		s_E902_C1_H				  :std_logic_vector(11 downto 0) := x"70C"; 
		s_E903_C1_H				  :std_logic_vector(11 downto 0) := x"70E"; 
		s_E904_C1_H				  :std_logic_vector(11 downto 0) := x"710"; 
		s_E905_C1_H				  :std_logic_vector(11 downto 0) := x"712"; 
		s_E906_C1_H				  :std_logic_vector(11 downto 0) := x"714"; 
		s_E907_C1_H				  :std_logic_vector(11 downto 0) := x"716"; 
		s_E908_C1_H				  :std_logic_vector(11 downto 0) := x"718"; 
		s_E909_C1_H				  :std_logic_vector(11 downto 0) := x"71A"; 
		s_E910_C1_H				  :std_logic_vector(11 downto 0) := x"71C"; 
		s_E911_C1_H				  :std_logic_vector(11 downto 0) := x"71E"; 
		s_E912_C1_H				  :std_logic_vector(11 downto 0) := x"720"; 
		s_E913_C1_H				  :std_logic_vector(11 downto 0) := x"722"; 
		s_E914_C1_H				  :std_logic_vector(11 downto 0) := x"724"; 
		s_E915_C1_H				  :std_logic_vector(11 downto 0) := x"726"; 
		s_E916_C1_H				  :std_logic_vector(11 downto 0) := x"728"; 
		s_E917_C1_H				  :std_logic_vector(11 downto 0) := x"72A"; 
		s_E918_C1_H				  :std_logic_vector(11 downto 0) := x"72C"; 
		s_E919_C1_H				  :std_logic_vector(11 downto 0) := x"72E"; 
		s_E920_C1_H				  :std_logic_vector(11 downto 0) := x"730"; 
		s_E921_C1_H				  :std_logic_vector(11 downto 0) := x"732"; 
		s_E922_C1_H				  :std_logic_vector(11 downto 0) := x"734"; 
		s_E923_C1_H				  :std_logic_vector(11 downto 0) := x"736"; 
		s_E924_C1_H				  :std_logic_vector(11 downto 0) := x"738"; 
		s_E925_C1_H				  :std_logic_vector(11 downto 0) := x"73A"; 
		s_E926_C1_H				  :std_logic_vector(11 downto 0) := x"73C"; 
		s_E927_C1_H				  :std_logic_vector(11 downto 0) := x"73E"; 
		s_E928_C1_H				  :std_logic_vector(11 downto 0) := x"740"; 
		s_E929_C1_H				  :std_logic_vector(11 downto 0) := x"742"; 
		s_E930_C1_H				  :std_logic_vector(11 downto 0) := x"744"; 
		s_E931_C1_H				  :std_logic_vector(11 downto 0) := x"746"; 
		s_E932_C1_H				  :std_logic_vector(11 downto 0) := x"748"; 
		s_E933_C1_H				  :std_logic_vector(11 downto 0) := x"74A"; 
		s_E934_C1_H				  :std_logic_vector(11 downto 0) := x"74C"; 
		s_E935_C1_H				  :std_logic_vector(11 downto 0) := x"74E"; 
		s_E936_C1_H				  :std_logic_vector(11 downto 0) := x"750"; 
		s_E937_C1_H				  :std_logic_vector(11 downto 0) := x"752"; 
		s_E938_C1_H				  :std_logic_vector(11 downto 0) := x"754"; 
		s_E939_C1_H				  :std_logic_vector(11 downto 0) := x"756"; 
		s_E940_C1_H				  :std_logic_vector(11 downto 0) := x"758"; 
		s_E941_C1_H				  :std_logic_vector(11 downto 0) := x"75A"; 
		s_E942_C1_H				  :std_logic_vector(11 downto 0) := x"75C"; 
		s_E943_C1_H				  :std_logic_vector(11 downto 0) := x"75E"; 
		s_E944_C1_H				  :std_logic_vector(11 downto 0) := x"760"; 
		s_E945_C1_H				  :std_logic_vector(11 downto 0) := x"762"; 
		s_E946_C1_H				  :std_logic_vector(11 downto 0) := x"764"; 
		s_E947_C1_H				  :std_logic_vector(11 downto 0) := x"766"; 
		s_E948_C1_H				  :std_logic_vector(11 downto 0) := x"768"; 
		s_E949_C1_H				  :std_logic_vector(11 downto 0) := x"76A"; 
		s_E950_C1_H				  :std_logic_vector(11 downto 0) := x"76C"; 
		s_E951_C1_H				  :std_logic_vector(11 downto 0) := x"76E"; 
		s_E952_C1_H				  :std_logic_vector(11 downto 0) := x"770"; 
		s_E953_C1_H				  :std_logic_vector(11 downto 0) := x"772"; 
		s_E954_C1_H				  :std_logic_vector(11 downto 0) := x"774"; 
		s_E955_C1_H				  :std_logic_vector(11 downto 0) := x"776"; 
		s_E956_C1_H				  :std_logic_vector(11 downto 0) := x"778"; 
		s_E957_C1_H				  :std_logic_vector(11 downto 0) := x"77A"; 
		s_E958_C1_H				  :std_logic_vector(11 downto 0) := x"77C"; 
		s_E959_C1_H				  :std_logic_vector(11 downto 0) := x"77E"; 
		s_E960_C1_H				  :std_logic_vector(11 downto 0) := x"780"; 
		s_E961_C1_H				  :std_logic_vector(11 downto 0) := x"782"; 
		s_E962_C1_H				  :std_logic_vector(11 downto 0) := x"784"; 
		s_E963_C1_H				  :std_logic_vector(11 downto 0) := x"786"; 
		s_E964_C1_H				  :std_logic_vector(11 downto 0) := x"788"; 
		s_E965_C1_H				  :std_logic_vector(11 downto 0) := x"78A"; 
		s_E966_C1_H				  :std_logic_vector(11 downto 0) := x"78C"; 
		s_E967_C1_H				  :std_logic_vector(11 downto 0) := x"78E"; 
		s_E968_C1_H				  :std_logic_vector(11 downto 0) := x"790"; 
		s_E969_C1_H				  :std_logic_vector(11 downto 0) := x"792"; 
		s_E970_C1_H				  :std_logic_vector(11 downto 0) := x"794"; 
		s_E971_C1_H				  :std_logic_vector(11 downto 0) := x"796"; 
		s_E972_C1_H				  :std_logic_vector(11 downto 0) := x"798"; 
		s_E973_C1_H				  :std_logic_vector(11 downto 0) := x"79A"; 
		s_E974_C1_H				  :std_logic_vector(11 downto 0) := x"79C"; 
		s_E975_C1_H				  :std_logic_vector(11 downto 0) := x"79E"; 
		s_E976_C1_H				  :std_logic_vector(11 downto 0) := x"7A0"; 
		s_E977_C1_H				  :std_logic_vector(11 downto 0) := x"7A2"; 
		s_E978_C1_H				  :std_logic_vector(11 downto 0) := x"7A4"; 
		s_E979_C1_H				  :std_logic_vector(11 downto 0) := x"7A6"; 
		s_E980_C1_H				  :std_logic_vector(11 downto 0) := x"7A8"; 
		s_E981_C1_H				  :std_logic_vector(11 downto 0) := x"7AA"; 
		s_E982_C1_H				  :std_logic_vector(11 downto 0) := x"7AC"; 
		s_E983_C1_H				  :std_logic_vector(11 downto 0) := x"7AE"; 
		s_E984_C1_H				  :std_logic_vector(11 downto 0) := x"7B0"; 
		s_E985_C1_H				  :std_logic_vector(11 downto 0) := x"7B2"; 
		s_E986_C1_H				  :std_logic_vector(11 downto 0) := x"7B4"; 
		s_E987_C1_H				  :std_logic_vector(11 downto 0) := x"7B6"; 
		s_E988_C1_H				  :std_logic_vector(11 downto 0) := x"7B8"; 
		s_E989_C1_H				  :std_logic_vector(11 downto 0) := x"7BA"; 
		s_E990_C1_H				  :std_logic_vector(11 downto 0) := x"7BC"; 
		s_E991_C1_H				  :std_logic_vector(11 downto 0) := x"7BE"; 
		s_E992_C1_H				  :std_logic_vector(11 downto 0) := x"7C0"; 
		s_E993_C1_H				  :std_logic_vector(11 downto 0) := x"7C2"; 
		s_E994_C1_H				  :std_logic_vector(11 downto 0) := x"7C4"; 
		s_E995_C1_H				  :std_logic_vector(11 downto 0) := x"7C6"; 
		s_E996_C1_H				  :std_logic_vector(11 downto 0) := x"7C8"; 
		s_E997_C1_H				  :std_logic_vector(11 downto 0) := x"7CA"; 
		s_E998_C1_H				  :std_logic_vector(11 downto 0) := x"7CC"; 
		s_E999_C1_H				  :std_logic_vector(11 downto 0) := x"7CE"; 
		s_E1000_C1_H			  :std_logic_vector(11 downto 0) := x"7D0"; 
		s_E1001_C1_H			  :std_logic_vector(11 downto 0) := x"7D2"; 
		s_E1002_C1_H			  :std_logic_vector(11 downto 0) := x"7D4"; 
		s_E1003_C1_H			  :std_logic_vector(11 downto 0) := x"7D6"; 
		s_E1004_C1_H			  :std_logic_vector(11 downto 0) := x"7D8"; 
		s_E1005_C1_H			  :std_logic_vector(11 downto 0) := x"7DA"; 
		s_E1006_C1_H			  :std_logic_vector(11 downto 0) := x"7DC"; 
		s_E1007_C1_H			  :std_logic_vector(11 downto 0) := x"7DE"; 
		s_E1008_C1_H			  :std_logic_vector(11 downto 0) := x"7E0"; 
		s_E1009_C1_H			  :std_logic_vector(11 downto 0) := x"7E2"; 
		s_E1010_C1_H			  :std_logic_vector(11 downto 0) := x"7E4"; 
		s_E1011_C1_H			  :std_logic_vector(11 downto 0) := x"7E6"; 
		s_E1012_C1_H			  :std_logic_vector(11 downto 0) := x"7E8"; 
		s_E1013_C1_H			  :std_logic_vector(11 downto 0) := x"7EA"; 
		s_E1014_C1_H			  :std_logic_vector(11 downto 0) := x"7EC"; 
		s_E1015_C1_H			  :std_logic_vector(11 downto 0) := x"7EE"; 
		s_E1016_C1_H			  :std_logic_vector(11 downto 0) := x"7F0"; 
		s_E1017_C1_H			  :std_logic_vector(11 downto 0) := x"7F2"; 
		s_E1018_C1_H			  :std_logic_vector(11 downto 0) := x"7F4"; 
		s_E1019_C1_H			  :std_logic_vector(11 downto 0) := x"7F6"; 
		s_E1020_C1_H			  :std_logic_vector(11 downto 0) := x"7F8"; 
		s_E1021_C1_H			  :std_logic_vector(11 downto 0) := x"7FA"; 
		s_E1022_C1_H			  :std_logic_vector(11 downto 0) := x"7FC"; 
		s_E1023_C1_H			  :std_logic_vector(11 downto 0) := x"7FE"; 
		s_E1024_C1_H			  :std_logic_vector(11 downto 0) := x"7FF"; 
		
		s_E2_C1_L       	 	  :std_logic_vector(11 downto 0) := x"002"; 
		s_E3_C1_L       	 	  :std_logic_vector(11 downto 0) := x"004"; 
		s_E4_C1_L       	 	  :std_logic_vector(11 downto 0) := x"006"; 
		s_E5_C1_L       	 	  :std_logic_vector(11 downto 0) := x"008"; 
		s_E6_C1_L       	 	  :std_logic_vector(11 downto 0) := x"00A"; 
		s_E7_C1_L       	 	  :std_logic_vector(11 downto 0) := x"00C"; 
		s_E8_C1_L       	 	  :std_logic_vector(11 downto 0) := x"00E"; 
		s_E9_C1_L       	 	  :std_logic_vector(11 downto 0) := x"010"; 
		s_E10_C1_L       	 	  :std_logic_vector(11 downto 0) := x"012"; 
		s_E11_C1_L				  :std_logic_vector(11 downto 0) := x"014"; 
		s_E12_C1_L				  :std_logic_vector(11 downto 0) := x"016"; 
		s_E13_C1_L				  :std_logic_vector(11 downto 0) := x"018"; 
		s_E14_C1_L				  :std_logic_vector(11 downto 0) := x"01A"; 
		s_E15_C1_L				  :std_logic_vector(11 downto 0) := x"01C"; 
		s_E16_C1_L				  :std_logic_vector(11 downto 0) := x"01E"; 
		s_E17_C1_L				  :std_logic_vector(11 downto 0) := x"020"; 
		s_E18_C1_L				  :std_logic_vector(11 downto 0) := x"022"; 
		s_E19_C1_L				  :std_logic_vector(11 downto 0) := x"024"; 
		s_E20_C1_L				  :std_logic_vector(11 downto 0) := x"026"; 
		s_E21_C1_L				  :std_logic_vector(11 downto 0) := x"028"; 
		s_E22_C1_L				  :std_logic_vector(11 downto 0) := x"02A"; 
		s_E23_C1_L				  :std_logic_vector(11 downto 0) := x"02C"; 
		s_E24_C1_L				  :std_logic_vector(11 downto 0) := x"02E"; 
		s_E25_C1_L				  :std_logic_vector(11 downto 0) := x"030"; 
		s_E26_C1_L				  :std_logic_vector(11 downto 0) := x"032"; 
		s_E27_C1_L				  :std_logic_vector(11 downto 0) := x"034"; 
		s_E28_C1_L				  :std_logic_vector(11 downto 0) := x"036"; 
		s_E29_C1_L				  :std_logic_vector(11 downto 0) := x"038"; 
		s_E30_C1_L				  :std_logic_vector(11 downto 0) := x"03A"; 
		s_E31_C1_L				  :std_logic_vector(11 downto 0) := x"03C"; 
		s_E32_C1_L				  :std_logic_vector(11 downto 0) := x"03E"; 
		s_E33_C1_L				  :std_logic_vector(11 downto 0) := x"040"; 
		s_E34_C1_L				  :std_logic_vector(11 downto 0) := x"042"; 
		s_E35_C1_L				  :std_logic_vector(11 downto 0) := x"044"; 
		s_E36_C1_L				  :std_logic_vector(11 downto 0) := x"046"; 
		s_E37_C1_L				  :std_logic_vector(11 downto 0) := x"048"; 
		s_E38_C1_L				  :std_logic_vector(11 downto 0) := x"04A"; 
		s_E39_C1_L				  :std_logic_vector(11 downto 0) := x"04C"; 
		s_E40_C1_L				  :std_logic_vector(11 downto 0) := x"04E"; 
		s_E41_C1_L				  :std_logic_vector(11 downto 0) := x"050"; 
		s_E42_C1_L				  :std_logic_vector(11 downto 0) := x"052"; 
		s_E43_C1_L				  :std_logic_vector(11 downto 0) := x"054"; 
		s_E44_C1_L				  :std_logic_vector(11 downto 0) := x"056"; 
		s_E45_C1_L				  :std_logic_vector(11 downto 0) := x"058"; 
		s_E46_C1_L				  :std_logic_vector(11 downto 0) := x"05A"; 
		s_E47_C1_L				  :std_logic_vector(11 downto 0) := x"05C"; 
		s_E48_C1_L				  :std_logic_vector(11 downto 0) := x"05E"; 
		s_E49_C1_L				  :std_logic_vector(11 downto 0) := x"060"; 
		s_E50_C1_L				  :std_logic_vector(11 downto 0) := x"062"; 
		s_E51_C1_L				  :std_logic_vector(11 downto 0) := x"064"; 
		s_E52_C1_L				  :std_logic_vector(11 downto 0) := x"066"; 
		s_E53_C1_L				  :std_logic_vector(11 downto 0) := x"068"; 
		s_E54_C1_L				  :std_logic_vector(11 downto 0) := x"06A"; 
		s_E55_C1_L				  :std_logic_vector(11 downto 0) := x"06C"; 
		s_E56_C1_L				  :std_logic_vector(11 downto 0) := x"06E"; 
		s_E57_C1_L				  :std_logic_vector(11 downto 0) := x"070"; 
		s_E58_C1_L				  :std_logic_vector(11 downto 0) := x"072"; 
		s_E59_C1_L				  :std_logic_vector(11 downto 0) := x"074"; 
		s_E60_C1_L				  :std_logic_vector(11 downto 0) := x"076"; 
		s_E61_C1_L				  :std_logic_vector(11 downto 0) := x"078"; 
		s_E62_C1_L				  :std_logic_vector(11 downto 0) := x"07A"; 
		s_E63_C1_L				  :std_logic_vector(11 downto 0) := x"07C"; 
		s_E64_C1_L				  :std_logic_vector(11 downto 0) := x"07E"; 
		s_E65_C1_L				  :std_logic_vector(11 downto 0) := x"080"; 
		s_E66_C1_L				  :std_logic_vector(11 downto 0) := x"082"; 
		s_E67_C1_L				  :std_logic_vector(11 downto 0) := x"084"; 
		s_E68_C1_L				  :std_logic_vector(11 downto 0) := x"086"; 
		s_E69_C1_L				  :std_logic_vector(11 downto 0) := x"088"; 
		s_E70_C1_L				  :std_logic_vector(11 downto 0) := x"08A"; 
		s_E71_C1_L				  :std_logic_vector(11 downto 0) := x"08C"; 
		s_E72_C1_L				  :std_logic_vector(11 downto 0) := x"08E"; 
		s_E73_C1_L				  :std_logic_vector(11 downto 0) := x"090"; 
		s_E74_C1_L				  :std_logic_vector(11 downto 0) := x"092"; 
		s_E75_C1_L				  :std_logic_vector(11 downto 0) := x"094"; 
		s_E76_C1_L				  :std_logic_vector(11 downto 0) := x"096"; 
		s_E77_C1_L				  :std_logic_vector(11 downto 0) := x"098"; 
		s_E78_C1_L				  :std_logic_vector(11 downto 0) := x"09A"; 
		s_E79_C1_L				  :std_logic_vector(11 downto 0) := x"09C"; 
		s_E80_C1_L				  :std_logic_vector(11 downto 0) := x"09E"; 
		s_E81_C1_L				  :std_logic_vector(11 downto 0) := x"0A0"; 
		s_E82_C1_L				  :std_logic_vector(11 downto 0) := x"0A2"; 
		s_E83_C1_L				  :std_logic_vector(11 downto 0) := x"0A4"; 
		s_E84_C1_L				  :std_logic_vector(11 downto 0) := x"0A6"; 
		s_E85_C1_L				  :std_logic_vector(11 downto 0) := x"0A8"; 
		s_E86_C1_L				  :std_logic_vector(11 downto 0) := x"0AA"; 
		s_E87_C1_L				  :std_logic_vector(11 downto 0) := x"0AC"; 
		s_E88_C1_L				  :std_logic_vector(11 downto 0) := x"0AE"; 
		s_E89_C1_L				  :std_logic_vector(11 downto 0) := x"0B0"; 
		s_E90_C1_L				  :std_logic_vector(11 downto 0) := x"0B2"; 
		s_E91_C1_L				  :std_logic_vector(11 downto 0) := x"0B4"; 
		s_E92_C1_L				  :std_logic_vector(11 downto 0) := x"0B6"; 
		s_E93_C1_L				  :std_logic_vector(11 downto 0) := x"0B8"; 
		s_E94_C1_L				  :std_logic_vector(11 downto 0) := x"0BA"; 
		s_E95_C1_L				  :std_logic_vector(11 downto 0) := x"0BC"; 
		s_E96_C1_L				  :std_logic_vector(11 downto 0) := x"0BE"; 
		s_E97_C1_L				  :std_logic_vector(11 downto 0) := x"0C0"; 
		s_E98_C1_L				  :std_logic_vector(11 downto 0) := x"0C2"; 
		s_E99_C1_L				  :std_logic_vector(11 downto 0) := x"0C4"; 
		s_E100_C1_L				  :std_logic_vector(11 downto 0) := x"0C6"; 
		s_E101_C1_L				  :std_logic_vector(11 downto 0) := x"0C8"; 
		s_E102_C1_L				  :std_logic_vector(11 downto 0) := x"0CA"; 
		s_E103_C1_L				  :std_logic_vector(11 downto 0) := x"0CC"; 
		s_E104_C1_L				  :std_logic_vector(11 downto 0) := x"0CE"; 
		s_E105_C1_L				  :std_logic_vector(11 downto 0) := x"0D0"; 
		s_E106_C1_L				  :std_logic_vector(11 downto 0) := x"0D2"; 
		s_E107_C1_L				  :std_logic_vector(11 downto 0) := x"0D4"; 
		s_E108_C1_L				  :std_logic_vector(11 downto 0) := x"0D6"; 
		s_E109_C1_L				  :std_logic_vector(11 downto 0) := x"0D8"; 
		s_E110_C1_L				  :std_logic_vector(11 downto 0) := x"0DA"; 
		s_E111_C1_L				  :std_logic_vector(11 downto 0) := x"0DC"; 
		s_E112_C1_L				  :std_logic_vector(11 downto 0) := x"0DE"; 
		s_E113_C1_L				  :std_logic_vector(11 downto 0) := x"0E0"; 
		s_E114_C1_L				  :std_logic_vector(11 downto 0) := x"0E2"; 
		s_E115_C1_L				  :std_logic_vector(11 downto 0) := x"0E4"; 
		s_E116_C1_L				  :std_logic_vector(11 downto 0) := x"0E6"; 
		s_E117_C1_L				  :std_logic_vector(11 downto 0) := x"0E8"; 
		s_E118_C1_L				  :std_logic_vector(11 downto 0) := x"0EA"; 
		s_E119_C1_L				  :std_logic_vector(11 downto 0) := x"0EC"; 
		s_E120_C1_L				  :std_logic_vector(11 downto 0) := x"0EE"; 
		s_E121_C1_L				  :std_logic_vector(11 downto 0) := x"0F0"; 
		s_E122_C1_L				  :std_logic_vector(11 downto 0) := x"0F2"; 
		s_E123_C1_L				  :std_logic_vector(11 downto 0) := x"0F4"; 
		s_E124_C1_L				  :std_logic_vector(11 downto 0) := x"0F6"; 
		s_E125_C1_L				  :std_logic_vector(11 downto 0) := x"0F8"; 
		s_E126_C1_L				  :std_logic_vector(11 downto 0) := x"0FA"; 
		s_E127_C1_L				  :std_logic_vector(11 downto 0) := x"0FC"; 
		s_E128_C1_L				  :std_logic_vector(11 downto 0) := x"0FE"; 
		s_E129_C1_L				  :std_logic_vector(11 downto 0) := x"100"; 
		s_E130_C1_L				  :std_logic_vector(11 downto 0) := x"102"; 
		s_E131_C1_L				  :std_logic_vector(11 downto 0) := x"104"; 
		s_E132_C1_L				  :std_logic_vector(11 downto 0) := x"106"; 
		s_E133_C1_L				  :std_logic_vector(11 downto 0) := x"108"; 
		s_E134_C1_L				  :std_logic_vector(11 downto 0) := x"10A"; 
		s_E135_C1_L				  :std_logic_vector(11 downto 0) := x"10C"; 
		s_E136_C1_L				  :std_logic_vector(11 downto 0) := x"10E"; 
		s_E137_C1_L				  :std_logic_vector(11 downto 0) := x"110"; 
		s_E138_C1_L				  :std_logic_vector(11 downto 0) := x"112"; 
		s_E139_C1_L				  :std_logic_vector(11 downto 0) := x"114"; 
		s_E140_C1_L				  :std_logic_vector(11 downto 0) := x"116"; 
		s_E141_C1_L				  :std_logic_vector(11 downto 0) := x"118"; 
		s_E142_C1_L				  :std_logic_vector(11 downto 0) := x"11A"; 
		s_E143_C1_L				  :std_logic_vector(11 downto 0) := x"11C"; 
		s_E144_C1_L				  :std_logic_vector(11 downto 0) := x"11E"; 
		s_E145_C1_L				  :std_logic_vector(11 downto 0) := x"120"; 
		s_E146_C1_L				  :std_logic_vector(11 downto 0) := x"122"; 
		s_E147_C1_L				  :std_logic_vector(11 downto 0) := x"124"; 
		s_E148_C1_L				  :std_logic_vector(11 downto 0) := x"126"; 
		s_E149_C1_L				  :std_logic_vector(11 downto 0) := x"128"; 
		s_E150_C1_L				  :std_logic_vector(11 downto 0) := x"12A"; 
		s_E151_C1_L				  :std_logic_vector(11 downto 0) := x"12C"; 
		s_E152_C1_L				  :std_logic_vector(11 downto 0) := x"12E"; 
		s_E153_C1_L				  :std_logic_vector(11 downto 0) := x"130"; 
		s_E154_C1_L				  :std_logic_vector(11 downto 0) := x"132"; 
		s_E155_C1_L				  :std_logic_vector(11 downto 0) := x"134"; 
		s_E156_C1_L				  :std_logic_vector(11 downto 0) := x"136"; 
		s_E157_C1_L				  :std_logic_vector(11 downto 0) := x"138"; 
		s_E158_C1_L				  :std_logic_vector(11 downto 0) := x"13A"; 
		s_E159_C1_L				  :std_logic_vector(11 downto 0) := x"13C"; 
		s_E160_C1_L				  :std_logic_vector(11 downto 0) := x"13E"; 
		s_E161_C1_L				  :std_logic_vector(11 downto 0) := x"140"; 
		s_E162_C1_L				  :std_logic_vector(11 downto 0) := x"142"; 
		s_E163_C1_L				  :std_logic_vector(11 downto 0) := x"144"; 
		s_E164_C1_L				  :std_logic_vector(11 downto 0) := x"146"; 
		s_E165_C1_L				  :std_logic_vector(11 downto 0) := x"148"; 
		s_E166_C1_L				  :std_logic_vector(11 downto 0) := x"14A"; 
		s_E167_C1_L				  :std_logic_vector(11 downto 0) := x"14C"; 
		s_E168_C1_L				  :std_logic_vector(11 downto 0) := x"14E"; 
		s_E169_C1_L				  :std_logic_vector(11 downto 0) := x"150"; 
		s_E170_C1_L				  :std_logic_vector(11 downto 0) := x"152"; 
		s_E171_C1_L				  :std_logic_vector(11 downto 0) := x"154"; 
		s_E172_C1_L				  :std_logic_vector(11 downto 0) := x"156"; 
		s_E173_C1_L				  :std_logic_vector(11 downto 0) := x"158"; 
		s_E174_C1_L				  :std_logic_vector(11 downto 0) := x"15A"; 
		s_E175_C1_L				  :std_logic_vector(11 downto 0) := x"15C"; 
		s_E176_C1_L				  :std_logic_vector(11 downto 0) := x"15E"; 
		s_E177_C1_L				  :std_logic_vector(11 downto 0) := x"160"; 
		s_E178_C1_L				  :std_logic_vector(11 downto 0) := x"162"; 
		s_E179_C1_L				  :std_logic_vector(11 downto 0) := x"164"; 
		s_E180_C1_L				  :std_logic_vector(11 downto 0) := x"166"; 
		s_E181_C1_L				  :std_logic_vector(11 downto 0) := x"168"; 
		s_E182_C1_L				  :std_logic_vector(11 downto 0) := x"16A"; 
		s_E183_C1_L				  :std_logic_vector(11 downto 0) := x"16C"; 
		s_E184_C1_L				  :std_logic_vector(11 downto 0) := x"16E"; 
		s_E185_C1_L				  :std_logic_vector(11 downto 0) := x"170"; 
		s_E186_C1_L				  :std_logic_vector(11 downto 0) := x"172"; 
		s_E187_C1_L				  :std_logic_vector(11 downto 0) := x"174"; 
		s_E188_C1_L				  :std_logic_vector(11 downto 0) := x"176"; 
		s_E189_C1_L				  :std_logic_vector(11 downto 0) := x"178"; 
		s_E190_C1_L				  :std_logic_vector(11 downto 0) := x"17A"; 
		s_E191_C1_L				  :std_logic_vector(11 downto 0) := x"17C"; 
		s_E192_C1_L				  :std_logic_vector(11 downto 0) := x"17E"; 
		s_E193_C1_L				  :std_logic_vector(11 downto 0) := x"180"; 
		s_E194_C1_L				  :std_logic_vector(11 downto 0) := x"182"; 
		s_E195_C1_L				  :std_logic_vector(11 downto 0) := x"184"; 
		s_E196_C1_L				  :std_logic_vector(11 downto 0) := x"186"; 
		s_E197_C1_L				  :std_logic_vector(11 downto 0) := x"188"; 
		s_E198_C1_L				  :std_logic_vector(11 downto 0) := x"18A"; 
		s_E199_C1_L				  :std_logic_vector(11 downto 0) := x"18C"; 
		s_E200_C1_L				  :std_logic_vector(11 downto 0) := x"18E"; 
		s_E201_C1_L				  :std_logic_vector(11 downto 0) := x"190"; 
		s_E202_C1_L				  :std_logic_vector(11 downto 0) := x"192"; 
		s_E203_C1_L				  :std_logic_vector(11 downto 0) := x"194"; 
		s_E204_C1_L				  :std_logic_vector(11 downto 0) := x"196"; 
		s_E205_C1_L				  :std_logic_vector(11 downto 0) := x"198"; 
		s_E206_C1_L				  :std_logic_vector(11 downto 0) := x"19A"; 
		s_E207_C1_L				  :std_logic_vector(11 downto 0) := x"19C"; 
		s_E208_C1_L				  :std_logic_vector(11 downto 0) := x"19E"; 
		s_E209_C1_L				  :std_logic_vector(11 downto 0) := x"1A0"; 
		s_E210_C1_L				  :std_logic_vector(11 downto 0) := x"1A2"; 
		s_E211_C1_L				  :std_logic_vector(11 downto 0) := x"1A4"; 
		s_E212_C1_L				  :std_logic_vector(11 downto 0) := x"1A6"; 
		s_E213_C1_L				  :std_logic_vector(11 downto 0) := x"1A8"; 
		s_E214_C1_L				  :std_logic_vector(11 downto 0) := x"1AA"; 
		s_E215_C1_L				  :std_logic_vector(11 downto 0) := x"1AC"; 
		s_E216_C1_L				  :std_logic_vector(11 downto 0) := x"1AE"; 
		s_E217_C1_L				  :std_logic_vector(11 downto 0) := x"1B0"; 
		s_E218_C1_L				  :std_logic_vector(11 downto 0) := x"1B2"; 
		s_E219_C1_L				  :std_logic_vector(11 downto 0) := x"1B4"; 
		s_E220_C1_L				  :std_logic_vector(11 downto 0) := x"1B6"; 
		s_E221_C1_L				  :std_logic_vector(11 downto 0) := x"1B8"; 
		s_E222_C1_L				  :std_logic_vector(11 downto 0) := x"1BA"; 
		s_E223_C1_L				  :std_logic_vector(11 downto 0) := x"1BC"; 
		s_E224_C1_L				  :std_logic_vector(11 downto 0) := x"1BE"; 
		s_E225_C1_L				  :std_logic_vector(11 downto 0) := x"1C0"; 
		s_E226_C1_L				  :std_logic_vector(11 downto 0) := x"1C2"; 
		s_E227_C1_L				  :std_logic_vector(11 downto 0) := x"1C4"; 
		s_E228_C1_L				  :std_logic_vector(11 downto 0) := x"1C6"; 
		s_E229_C1_L				  :std_logic_vector(11 downto 0) := x"1C8"; 
		s_E230_C1_L				  :std_logic_vector(11 downto 0) := x"1CA"; 
		s_E231_C1_L				  :std_logic_vector(11 downto 0) := x"1CC"; 
		s_E232_C1_L				  :std_logic_vector(11 downto 0) := x"1CE"; 
		s_E233_C1_L				  :std_logic_vector(11 downto 0) := x"1D0"; 
		s_E234_C1_L				  :std_logic_vector(11 downto 0) := x"1D2"; 
		s_E235_C1_L				  :std_logic_vector(11 downto 0) := x"1D4"; 
		s_E236_C1_L				  :std_logic_vector(11 downto 0) := x"1D6"; 
		s_E237_C1_L				  :std_logic_vector(11 downto 0) := x"1D8"; 
		s_E238_C1_L				  :std_logic_vector(11 downto 0) := x"1DA"; 
		s_E239_C1_L				  :std_logic_vector(11 downto 0) := x"1DC"; 
		s_E240_C1_L				  :std_logic_vector(11 downto 0) := x"1DE"; 
		s_E241_C1_L				  :std_logic_vector(11 downto 0) := x"1E0"; 
		s_E242_C1_L				  :std_logic_vector(11 downto 0) := x"1E2"; 
		s_E243_C1_L				  :std_logic_vector(11 downto 0) := x"1E4"; 
		s_E244_C1_L				  :std_logic_vector(11 downto 0) := x"1E6"; 
		s_E245_C1_L				  :std_logic_vector(11 downto 0) := x"1E8"; 
		s_E246_C1_L				  :std_logic_vector(11 downto 0) := x"1EA"; 
		s_E247_C1_L				  :std_logic_vector(11 downto 0) := x"1EC"; 
		s_E248_C1_L				  :std_logic_vector(11 downto 0) := x"1EE"; 
		s_E249_C1_L				  :std_logic_vector(11 downto 0) := x"1F0"; 
		s_E250_C1_L				  :std_logic_vector(11 downto 0) := x"1F2"; 
		s_E251_C1_L				  :std_logic_vector(11 downto 0) := x"1F4"; 
		s_E252_C1_L				  :std_logic_vector(11 downto 0) := x"1F6"; 
		s_E253_C1_L				  :std_logic_vector(11 downto 0) := x"1F8"; 
		s_E254_C1_L				  :std_logic_vector(11 downto 0) := x"1FA"; 
		s_E255_C1_L				  :std_logic_vector(11 downto 0) := x"1FC"; 
		s_E256_C1_L				  :std_logic_vector(11 downto 0) := x"1FE"; 
		s_E257_C1_L				  :std_logic_vector(11 downto 0) := x"200"; 
		s_E258_C1_L				  :std_logic_vector(11 downto 0) := x"202"; 
		s_E259_C1_L				  :std_logic_vector(11 downto 0) := x"204"; 
		s_E260_C1_L				  :std_logic_vector(11 downto 0) := x"206"; 
		s_E261_C1_L				  :std_logic_vector(11 downto 0) := x"208"; 
		s_E262_C1_L				  :std_logic_vector(11 downto 0) := x"20A"; 
		s_E263_C1_L				  :std_logic_vector(11 downto 0) := x"20C"; 
		s_E264_C1_L				  :std_logic_vector(11 downto 0) := x"20E"; 
		s_E265_C1_L				  :std_logic_vector(11 downto 0) := x"210"; 
		s_E266_C1_L				  :std_logic_vector(11 downto 0) := x"212"; 
		s_E267_C1_L				  :std_logic_vector(11 downto 0) := x"214"; 
		s_E268_C1_L				  :std_logic_vector(11 downto 0) := x"216"; 
		s_E269_C1_L				  :std_logic_vector(11 downto 0) := x"218"; 
		s_E270_C1_L				  :std_logic_vector(11 downto 0) := x"21A"; 
		s_E271_C1_L				  :std_logic_vector(11 downto 0) := x"21C"; 
		s_E272_C1_L				  :std_logic_vector(11 downto 0) := x"21E"; 
		s_E273_C1_L				  :std_logic_vector(11 downto 0) := x"220"; 
		s_E274_C1_L				  :std_logic_vector(11 downto 0) := x"222"; 
		s_E275_C1_L				  :std_logic_vector(11 downto 0) := x"224"; 
		s_E276_C1_L				  :std_logic_vector(11 downto 0) := x"226"; 
		s_E277_C1_L				  :std_logic_vector(11 downto 0) := x"228"; 
		s_E278_C1_L				  :std_logic_vector(11 downto 0) := x"22A"; 
		s_E279_C1_L				  :std_logic_vector(11 downto 0) := x"22C"; 
		s_E280_C1_L				  :std_logic_vector(11 downto 0) := x"22E"; 
		s_E281_C1_L				  :std_logic_vector(11 downto 0) := x"230"; 
		s_E282_C1_L				  :std_logic_vector(11 downto 0) := x"232"; 
		s_E283_C1_L				  :std_logic_vector(11 downto 0) := x"234"; 
		s_E284_C1_L				  :std_logic_vector(11 downto 0) := x"236"; 
		s_E285_C1_L				  :std_logic_vector(11 downto 0) := x"238"; 
		s_E286_C1_L				  :std_logic_vector(11 downto 0) := x"23A"; 
		s_E287_C1_L				  :std_logic_vector(11 downto 0) := x"23C"; 
		s_E288_C1_L				  :std_logic_vector(11 downto 0) := x"23E"; 
		s_E289_C1_L				  :std_logic_vector(11 downto 0) := x"240"; 
		s_E290_C1_L				  :std_logic_vector(11 downto 0) := x"242"; 
		s_E291_C1_L				  :std_logic_vector(11 downto 0) := x"244"; 
		s_E292_C1_L				  :std_logic_vector(11 downto 0) := x"246"; 
		s_E293_C1_L				  :std_logic_vector(11 downto 0) := x"248"; 
		s_E294_C1_L				  :std_logic_vector(11 downto 0) := x"24A"; 
		s_E295_C1_L				  :std_logic_vector(11 downto 0) := x"24C"; 
		s_E296_C1_L				  :std_logic_vector(11 downto 0) := x"24E"; 
		s_E297_C1_L				  :std_logic_vector(11 downto 0) := x"250"; 
		s_E298_C1_L				  :std_logic_vector(11 downto 0) := x"252"; 
		s_E299_C1_L				  :std_logic_vector(11 downto 0) := x"254"; 
		s_E300_C1_L				  :std_logic_vector(11 downto 0) := x"256"; 
		s_E301_C1_L				  :std_logic_vector(11 downto 0) := x"258"; 
		s_E302_C1_L				  :std_logic_vector(11 downto 0) := x"25A"; 
		s_E303_C1_L				  :std_logic_vector(11 downto 0) := x"25C"; 
		s_E304_C1_L				  :std_logic_vector(11 downto 0) := x"25E"; 
		s_E305_C1_L				  :std_logic_vector(11 downto 0) := x"260"; 
		s_E306_C1_L				  :std_logic_vector(11 downto 0) := x"262"; 
		s_E307_C1_L				  :std_logic_vector(11 downto 0) := x"264"; 
		s_E308_C1_L				  :std_logic_vector(11 downto 0) := x"266"; 
		s_E309_C1_L				  :std_logic_vector(11 downto 0) := x"268"; 
		s_E310_C1_L				  :std_logic_vector(11 downto 0) := x"26A"; 
		s_E311_C1_L				  :std_logic_vector(11 downto 0) := x"26C"; 
		s_E312_C1_L				  :std_logic_vector(11 downto 0) := x"26E"; 
		s_E313_C1_L				  :std_logic_vector(11 downto 0) := x"270"; 
		s_E314_C1_L				  :std_logic_vector(11 downto 0) := x"272"; 
		s_E315_C1_L				  :std_logic_vector(11 downto 0) := x"274"; 
		s_E316_C1_L				  :std_logic_vector(11 downto 0) := x"276"; 
		s_E317_C1_L				  :std_logic_vector(11 downto 0) := x"278"; 
		s_E318_C1_L				  :std_logic_vector(11 downto 0) := x"27A"; 
		s_E319_C1_L				  :std_logic_vector(11 downto 0) := x"27C"; 
		s_E320_C1_L				  :std_logic_vector(11 downto 0) := x"27E"; 
		s_E321_C1_L				  :std_logic_vector(11 downto 0) := x"280"; 
		s_E322_C1_L				  :std_logic_vector(11 downto 0) := x"282"; 
		s_E323_C1_L				  :std_logic_vector(11 downto 0) := x"284"; 
		s_E324_C1_L				  :std_logic_vector(11 downto 0) := x"286"; 
		s_E325_C1_L				  :std_logic_vector(11 downto 0) := x"288"; 
		s_E326_C1_L				  :std_logic_vector(11 downto 0) := x"28A"; 
		s_E327_C1_L				  :std_logic_vector(11 downto 0) := x"28C"; 
		s_E328_C1_L				  :std_logic_vector(11 downto 0) := x"28E"; 
		s_E329_C1_L				  :std_logic_vector(11 downto 0) := x"290"; 
		s_E330_C1_L				  :std_logic_vector(11 downto 0) := x"292"; 
		s_E331_C1_L				  :std_logic_vector(11 downto 0) := x"294"; 
		s_E332_C1_L				  :std_logic_vector(11 downto 0) := x"296"; 
		s_E333_C1_L				  :std_logic_vector(11 downto 0) := x"298"; 
		s_E334_C1_L				  :std_logic_vector(11 downto 0) := x"29A"; 
		s_E335_C1_L				  :std_logic_vector(11 downto 0) := x"29C"; 
		s_E336_C1_L				  :std_logic_vector(11 downto 0) := x"29E"; 
		s_E337_C1_L				  :std_logic_vector(11 downto 0) := x"2A0"; 
		s_E338_C1_L				  :std_logic_vector(11 downto 0) := x"2A2"; 
		s_E339_C1_L				  :std_logic_vector(11 downto 0) := x"2A4"; 
		s_E340_C1_L				  :std_logic_vector(11 downto 0) := x"2A6"; 
		s_E341_C1_L				  :std_logic_vector(11 downto 0) := x"2A8"; 
		s_E342_C1_L				  :std_logic_vector(11 downto 0) := x"2AA"; 
		s_E343_C1_L				  :std_logic_vector(11 downto 0) := x"2AC"; 
		s_E344_C1_L				  :std_logic_vector(11 downto 0) := x"2AE"; 
		s_E345_C1_L				  :std_logic_vector(11 downto 0) := x"2B0"; 
		s_E346_C1_L				  :std_logic_vector(11 downto 0) := x"2B2"; 
		s_E347_C1_L				  :std_logic_vector(11 downto 0) := x"2B4"; 
		s_E348_C1_L				  :std_logic_vector(11 downto 0) := x"2B6"; 
		s_E349_C1_L				  :std_logic_vector(11 downto 0) := x"2B8"; 
		s_E350_C1_L				  :std_logic_vector(11 downto 0) := x"2BA"; 
		s_E351_C1_L				  :std_logic_vector(11 downto 0) := x"2BC"; 
		s_E352_C1_L				  :std_logic_vector(11 downto 0) := x"2BE"; 
		s_E353_C1_L				  :std_logic_vector(11 downto 0) := x"2C0"; 
		s_E354_C1_L				  :std_logic_vector(11 downto 0) := x"2C2"; 
		s_E355_C1_L				  :std_logic_vector(11 downto 0) := x"2C4"; 
		s_E356_C1_L				  :std_logic_vector(11 downto 0) := x"2C6"; 
		s_E357_C1_L				  :std_logic_vector(11 downto 0) := x"2C8"; 
		s_E358_C1_L				  :std_logic_vector(11 downto 0) := x"2CA"; 
		s_E359_C1_L				  :std_logic_vector(11 downto 0) := x"2CC"; 
		s_E360_C1_L				  :std_logic_vector(11 downto 0) := x"2CE"; 
		s_E361_C1_L				  :std_logic_vector(11 downto 0) := x"2D0"; 
		s_E362_C1_L				  :std_logic_vector(11 downto 0) := x"2D2"; 
		s_E363_C1_L				  :std_logic_vector(11 downto 0) := x"2D4"; 
		s_E364_C1_L				  :std_logic_vector(11 downto 0) := x"2D6"; 
		s_E365_C1_L				  :std_logic_vector(11 downto 0) := x"2D8"; 
		s_E366_C1_L				  :std_logic_vector(11 downto 0) := x"2DA"; 
		s_E367_C1_L				  :std_logic_vector(11 downto 0) := x"2DC"; 
		s_E368_C1_L				  :std_logic_vector(11 downto 0) := x"2DE"; 
		s_E369_C1_L				  :std_logic_vector(11 downto 0) := x"2E0"; 
		s_E370_C1_L				  :std_logic_vector(11 downto 0) := x"2E2"; 
		s_E371_C1_L				  :std_logic_vector(11 downto 0) := x"2E4"; 
		s_E372_C1_L				  :std_logic_vector(11 downto 0) := x"2E6"; 
		s_E373_C1_L				  :std_logic_vector(11 downto 0) := x"2E8"; 
		s_E374_C1_L				  :std_logic_vector(11 downto 0) := x"2EA"; 
		s_E375_C1_L				  :std_logic_vector(11 downto 0) := x"2EC"; 
		s_E376_C1_L				  :std_logic_vector(11 downto 0) := x"2EE"; 
		s_E377_C1_L				  :std_logic_vector(11 downto 0) := x"2F0"; 
		s_E378_C1_L				  :std_logic_vector(11 downto 0) := x"2F2"; 
		s_E379_C1_L				  :std_logic_vector(11 downto 0) := x"2F4"; 
		s_E380_C1_L				  :std_logic_vector(11 downto 0) := x"2F6"; 
		s_E381_C1_L				  :std_logic_vector(11 downto 0) := x"2F8"; 
		s_E382_C1_L				  :std_logic_vector(11 downto 0) := x"2FA"; 
		s_E383_C1_L				  :std_logic_vector(11 downto 0) := x"2FC"; 
		s_E384_C1_L				  :std_logic_vector(11 downto 0) := x"2FE"; 
		s_E385_C1_L				  :std_logic_vector(11 downto 0) := x"300"; 
		s_E386_C1_L				  :std_logic_vector(11 downto 0) := x"302"; 
		s_E387_C1_L				  :std_logic_vector(11 downto 0) := x"304"; 
		s_E388_C1_L				  :std_logic_vector(11 downto 0) := x"306"; 
		s_E389_C1_L				  :std_logic_vector(11 downto 0) := x"308"; 
		s_E390_C1_L				  :std_logic_vector(11 downto 0) := x"30A"; 
		s_E391_C1_L				  :std_logic_vector(11 downto 0) := x"30C"; 
		s_E392_C1_L				  :std_logic_vector(11 downto 0) := x"30E"; 
		s_E393_C1_L				  :std_logic_vector(11 downto 0) := x"310"; 
		s_E394_C1_L				  :std_logic_vector(11 downto 0) := x"312"; 
		s_E395_C1_L				  :std_logic_vector(11 downto 0) := x"314"; 
		s_E396_C1_L				  :std_logic_vector(11 downto 0) := x"316"; 
		s_E397_C1_L				  :std_logic_vector(11 downto 0) := x"318"; 
		s_E398_C1_L				  :std_logic_vector(11 downto 0) := x"31A"; 
		s_E399_C1_L				  :std_logic_vector(11 downto 0) := x"31C"; 
		s_E400_C1_L				  :std_logic_vector(11 downto 0) := x"31E"; 
		s_E401_C1_L				  :std_logic_vector(11 downto 0) := x"320"; 
		s_E402_C1_L				  :std_logic_vector(11 downto 0) := x"322"; 
		s_E403_C1_L				  :std_logic_vector(11 downto 0) := x"324"; 
		s_E404_C1_L				  :std_logic_vector(11 downto 0) := x"326"; 
		s_E405_C1_L				  :std_logic_vector(11 downto 0) := x"328"; 
		s_E406_C1_L				  :std_logic_vector(11 downto 0) := x"32A"; 
		s_E407_C1_L				  :std_logic_vector(11 downto 0) := x"32C"; 
		s_E408_C1_L				  :std_logic_vector(11 downto 0) := x"32E"; 
		s_E409_C1_L				  :std_logic_vector(11 downto 0) := x"330"; 
		s_E410_C1_L				  :std_logic_vector(11 downto 0) := x"332"; 
		s_E411_C1_L				  :std_logic_vector(11 downto 0) := x"334"; 
		s_E412_C1_L				  :std_logic_vector(11 downto 0) := x"336"; 
		s_E413_C1_L				  :std_logic_vector(11 downto 0) := x"338"; 
		s_E414_C1_L				  :std_logic_vector(11 downto 0) := x"33A"; 
		s_E415_C1_L				  :std_logic_vector(11 downto 0) := x"33C"; 
		s_E416_C1_L				  :std_logic_vector(11 downto 0) := x"33E"; 
		s_E417_C1_L				  :std_logic_vector(11 downto 0) := x"340"; 
		s_E418_C1_L				  :std_logic_vector(11 downto 0) := x"342"; 
		s_E419_C1_L				  :std_logic_vector(11 downto 0) := x"344"; 
		s_E420_C1_L				  :std_logic_vector(11 downto 0) := x"346"; 
		s_E421_C1_L				  :std_logic_vector(11 downto 0) := x"348"; 
		s_E422_C1_L				  :std_logic_vector(11 downto 0) := x"34A"; 
		s_E423_C1_L				  :std_logic_vector(11 downto 0) := x"34C"; 
		s_E424_C1_L				  :std_logic_vector(11 downto 0) := x"34E"; 
		s_E425_C1_L				  :std_logic_vector(11 downto 0) := x"350"; 
		s_E426_C1_L				  :std_logic_vector(11 downto 0) := x"352"; 
		s_E427_C1_L				  :std_logic_vector(11 downto 0) := x"354"; 
		s_E428_C1_L				  :std_logic_vector(11 downto 0) := x"356"; 
		s_E429_C1_L				  :std_logic_vector(11 downto 0) := x"358"; 
		s_E430_C1_L				  :std_logic_vector(11 downto 0) := x"35A"; 
		s_E431_C1_L				  :std_logic_vector(11 downto 0) := x"35C"; 
		s_E432_C1_L				  :std_logic_vector(11 downto 0) := x"35E"; 
		s_E433_C1_L				  :std_logic_vector(11 downto 0) := x"360"; 
		s_E434_C1_L				  :std_logic_vector(11 downto 0) := x"362"; 
		s_E435_C1_L				  :std_logic_vector(11 downto 0) := x"364"; 
		s_E436_C1_L				  :std_logic_vector(11 downto 0) := x"366"; 
		s_E437_C1_L				  :std_logic_vector(11 downto 0) := x"368"; 
		s_E438_C1_L				  :std_logic_vector(11 downto 0) := x"36A"; 
		s_E439_C1_L				  :std_logic_vector(11 downto 0) := x"36C"; 
		s_E440_C1_L				  :std_logic_vector(11 downto 0) := x"36E"; 
		s_E441_C1_L				  :std_logic_vector(11 downto 0) := x"370"; 
		s_E442_C1_L				  :std_logic_vector(11 downto 0) := x"372"; 
		s_E443_C1_L				  :std_logic_vector(11 downto 0) := x"374"; 
		s_E444_C1_L				  :std_logic_vector(11 downto 0) := x"376"; 
		s_E445_C1_L				  :std_logic_vector(11 downto 0) := x"378"; 
		s_E446_C1_L				  :std_logic_vector(11 downto 0) := x"37A"; 
		s_E447_C1_L				  :std_logic_vector(11 downto 0) := x"37C"; 
		s_E448_C1_L				  :std_logic_vector(11 downto 0) := x"37E"; 
		s_E449_C1_L				  :std_logic_vector(11 downto 0) := x"380"; 
		s_E450_C1_L				  :std_logic_vector(11 downto 0) := x"382"; 
		s_E451_C1_L				  :std_logic_vector(11 downto 0) := x"384"; 
		s_E452_C1_L				  :std_logic_vector(11 downto 0) := x"386"; 
		s_E453_C1_L				  :std_logic_vector(11 downto 0) := x"388"; 
		s_E454_C1_L				  :std_logic_vector(11 downto 0) := x"38A"; 
		s_E455_C1_L				  :std_logic_vector(11 downto 0) := x"38C"; 
		s_E456_C1_L				  :std_logic_vector(11 downto 0) := x"38E"; 
		s_E457_C1_L				  :std_logic_vector(11 downto 0) := x"390"; 
		s_E458_C1_L				  :std_logic_vector(11 downto 0) := x"392"; 
		s_E459_C1_L				  :std_logic_vector(11 downto 0) := x"394"; 
		s_E460_C1_L				  :std_logic_vector(11 downto 0) := x"396"; 
		s_E461_C1_L				  :std_logic_vector(11 downto 0) := x"398"; 
		s_E462_C1_L				  :std_logic_vector(11 downto 0) := x"39A"; 
		s_E463_C1_L				  :std_logic_vector(11 downto 0) := x"39C"; 
		s_E464_C1_L				  :std_logic_vector(11 downto 0) := x"39E"; 
		s_E465_C1_L				  :std_logic_vector(11 downto 0) := x"3A0"; 
		s_E466_C1_L				  :std_logic_vector(11 downto 0) := x"3A2"; 
		s_E467_C1_L				  :std_logic_vector(11 downto 0) := x"3A4"; 
		s_E468_C1_L				  :std_logic_vector(11 downto 0) := x"3A6"; 
		s_E469_C1_L				  :std_logic_vector(11 downto 0) := x"3A8"; 
		s_E470_C1_L				  :std_logic_vector(11 downto 0) := x"3AA"; 
		s_E471_C1_L				  :std_logic_vector(11 downto 0) := x"3AC"; 
		s_E472_C1_L				  :std_logic_vector(11 downto 0) := x"3AE"; 
		s_E473_C1_L				  :std_logic_vector(11 downto 0) := x"3B0"; 
		s_E474_C1_L				  :std_logic_vector(11 downto 0) := x"3B2"; 
		s_E475_C1_L				  :std_logic_vector(11 downto 0) := x"3B4"; 
		s_E476_C1_L				  :std_logic_vector(11 downto 0) := x"3B6"; 
		s_E477_C1_L				  :std_logic_vector(11 downto 0) := x"3B8"; 
		s_E478_C1_L				  :std_logic_vector(11 downto 0) := x"3BA"; 
		s_E479_C1_L				  :std_logic_vector(11 downto 0) := x"3BC"; 
		s_E480_C1_L				  :std_logic_vector(11 downto 0) := x"3BE"; 
		s_E481_C1_L				  :std_logic_vector(11 downto 0) := x"3C0"; 
		s_E482_C1_L				  :std_logic_vector(11 downto 0) := x"3C2"; 
		s_E483_C1_L				  :std_logic_vector(11 downto 0) := x"3C4"; 
		s_E484_C1_L				  :std_logic_vector(11 downto 0) := x"3C6"; 
		s_E485_C1_L				  :std_logic_vector(11 downto 0) := x"3C8"; 
		s_E486_C1_L				  :std_logic_vector(11 downto 0) := x"3CA"; 
		s_E487_C1_L				  :std_logic_vector(11 downto 0) := x"3CC"; 
		s_E488_C1_L				  :std_logic_vector(11 downto 0) := x"3CE"; 
		s_E489_C1_L				  :std_logic_vector(11 downto 0) := x"3D0"; 
		s_E490_C1_L				  :std_logic_vector(11 downto 0) := x"3D2"; 
		s_E491_C1_L				  :std_logic_vector(11 downto 0) := x"3D4"; 
		s_E492_C1_L				  :std_logic_vector(11 downto 0) := x"3D6"; 
		s_E493_C1_L				  :std_logic_vector(11 downto 0) := x"3D8"; 
		s_E494_C1_L				  :std_logic_vector(11 downto 0) := x"3DA"; 
		s_E495_C1_L				  :std_logic_vector(11 downto 0) := x"3DC"; 
		s_E496_C1_L				  :std_logic_vector(11 downto 0) := x"3DE"; 
		s_E497_C1_L				  :std_logic_vector(11 downto 0) := x"3E0"; 
		s_E498_C1_L				  :std_logic_vector(11 downto 0) := x"3E2"; 
		s_E499_C1_L				  :std_logic_vector(11 downto 0) := x"3E4"; 
		s_E500_C1_L				  :std_logic_vector(11 downto 0) := x"3E6"; 
		s_E501_C1_L				  :std_logic_vector(11 downto 0) := x"3E8"; 
		s_E502_C1_L				  :std_logic_vector(11 downto 0) := x"3EA"; 
		s_E503_C1_L				  :std_logic_vector(11 downto 0) := x"3EC"; 
		s_E504_C1_L				  :std_logic_vector(11 downto 0) := x"3EE"; 
		s_E505_C1_L				  :std_logic_vector(11 downto 0) := x"3F0"; 
		s_E506_C1_L				  :std_logic_vector(11 downto 0) := x"3F2"; 
		s_E507_C1_L				  :std_logic_vector(11 downto 0) := x"3F4"; 
		s_E508_C1_L				  :std_logic_vector(11 downto 0) := x"3F6"; 
		s_E509_C1_L				  :std_logic_vector(11 downto 0) := x"3F8"; 
		s_E510_C1_L				  :std_logic_vector(11 downto 0) := x"3FA"; 
		s_E511_C1_L				  :std_logic_vector(11 downto 0) := x"3FC"; 
		s_E512_C1_L				  :std_logic_vector(11 downto 0) := x"3FE"; 
		s_E513_C1_L				  :std_logic_vector(11 downto 0) := x"400"; 
		s_E514_C1_L				  :std_logic_vector(11 downto 0) := x"402"; 
		s_E515_C1_L				  :std_logic_vector(11 downto 0) := x"404"; 
		s_E516_C1_L				  :std_logic_vector(11 downto 0) := x"406"; 
		s_E517_C1_L				  :std_logic_vector(11 downto 0) := x"408"; 
		s_E518_C1_L				  :std_logic_vector(11 downto 0) := x"40A"; 
		s_E519_C1_L				  :std_logic_vector(11 downto 0) := x"40C"; 
		s_E520_C1_L				  :std_logic_vector(11 downto 0) := x"40E"; 
		s_E521_C1_L				  :std_logic_vector(11 downto 0) := x"410"; 
		s_E522_C1_L				  :std_logic_vector(11 downto 0) := x"412"; 
		s_E523_C1_L				  :std_logic_vector(11 downto 0) := x"414"; 
		s_E524_C1_L				  :std_logic_vector(11 downto 0) := x"416"; 
		s_E525_C1_L				  :std_logic_vector(11 downto 0) := x"418"; 
		s_E526_C1_L				  :std_logic_vector(11 downto 0) := x"41A"; 
		s_E527_C1_L				  :std_logic_vector(11 downto 0) := x"41C"; 
		s_E528_C1_L				  :std_logic_vector(11 downto 0) := x"41E"; 
		s_E529_C1_L				  :std_logic_vector(11 downto 0) := x"420"; 
		s_E530_C1_L				  :std_logic_vector(11 downto 0) := x"422"; 
		s_E531_C1_L				  :std_logic_vector(11 downto 0) := x"424"; 
		s_E532_C1_L				  :std_logic_vector(11 downto 0) := x"426"; 
		s_E533_C1_L				  :std_logic_vector(11 downto 0) := x"428"; 
		s_E534_C1_L				  :std_logic_vector(11 downto 0) := x"42A"; 
		s_E535_C1_L				  :std_logic_vector(11 downto 0) := x"42C"; 
		s_E536_C1_L				  :std_logic_vector(11 downto 0) := x"42E"; 
		s_E537_C1_L				  :std_logic_vector(11 downto 0) := x"430"; 
		s_E538_C1_L				  :std_logic_vector(11 downto 0) := x"432"; 
		s_E539_C1_L				  :std_logic_vector(11 downto 0) := x"434"; 
		s_E540_C1_L				  :std_logic_vector(11 downto 0) := x"436"; 
		s_E541_C1_L				  :std_logic_vector(11 downto 0) := x"438"; 
		s_E542_C1_L				  :std_logic_vector(11 downto 0) := x"43A"; 
		s_E543_C1_L				  :std_logic_vector(11 downto 0) := x"43C"; 
		s_E544_C1_L				  :std_logic_vector(11 downto 0) := x"43E"; 
		s_E545_C1_L				  :std_logic_vector(11 downto 0) := x"440"; 
		s_E546_C1_L				  :std_logic_vector(11 downto 0) := x"442"; 
		s_E547_C1_L				  :std_logic_vector(11 downto 0) := x"444"; 
		s_E548_C1_L				  :std_logic_vector(11 downto 0) := x"446"; 
		s_E549_C1_L				  :std_logic_vector(11 downto 0) := x"448"; 
		s_E550_C1_L				  :std_logic_vector(11 downto 0) := x"44A"; 
		s_E551_C1_L				  :std_logic_vector(11 downto 0) := x"44C"; 
		s_E552_C1_L				  :std_logic_vector(11 downto 0) := x"44E"; 
		s_E553_C1_L				  :std_logic_vector(11 downto 0) := x"450"; 
		s_E554_C1_L				  :std_logic_vector(11 downto 0) := x"452"; 
		s_E555_C1_L				  :std_logic_vector(11 downto 0) := x"454"; 
		s_E556_C1_L				  :std_logic_vector(11 downto 0) := x"456"; 
		s_E557_C1_L				  :std_logic_vector(11 downto 0) := x"458"; 
		s_E558_C1_L				  :std_logic_vector(11 downto 0) := x"45A"; 
		s_E559_C1_L				  :std_logic_vector(11 downto 0) := x"45C"; 
		s_E560_C1_L				  :std_logic_vector(11 downto 0) := x"45E"; 
		s_E561_C1_L				  :std_logic_vector(11 downto 0) := x"460"; 
		s_E562_C1_L				  :std_logic_vector(11 downto 0) := x"462"; 
		s_E563_C1_L				  :std_logic_vector(11 downto 0) := x"464"; 
		s_E564_C1_L				  :std_logic_vector(11 downto 0) := x"466"; 
		s_E565_C1_L				  :std_logic_vector(11 downto 0) := x"468"; 
		s_E566_C1_L				  :std_logic_vector(11 downto 0) := x"46A"; 
		s_E567_C1_L				  :std_logic_vector(11 downto 0) := x"46C"; 
		s_E568_C1_L				  :std_logic_vector(11 downto 0) := x"46E"; 
		s_E569_C1_L				  :std_logic_vector(11 downto 0) := x"470"; 
		s_E570_C1_L				  :std_logic_vector(11 downto 0) := x"472"; 
		s_E571_C1_L				  :std_logic_vector(11 downto 0) := x"474"; 
		s_E572_C1_L				  :std_logic_vector(11 downto 0) := x"476"; 
		s_E573_C1_L				  :std_logic_vector(11 downto 0) := x"478"; 
		s_E574_C1_L				  :std_logic_vector(11 downto 0) := x"47A"; 
		s_E575_C1_L				  :std_logic_vector(11 downto 0) := x"47C"; 
		s_E576_C1_L				  :std_logic_vector(11 downto 0) := x"47E"; 
		s_E577_C1_L				  :std_logic_vector(11 downto 0) := x"480"; 
		s_E578_C1_L				  :std_logic_vector(11 downto 0) := x"482"; 
		s_E579_C1_L				  :std_logic_vector(11 downto 0) := x"484"; 
		s_E580_C1_L				  :std_logic_vector(11 downto 0) := x"486"; 
		s_E581_C1_L				  :std_logic_vector(11 downto 0) := x"488"; 
		s_E582_C1_L				  :std_logic_vector(11 downto 0) := x"48A"; 
		s_E583_C1_L				  :std_logic_vector(11 downto 0) := x"48C"; 
		s_E584_C1_L				  :std_logic_vector(11 downto 0) := x"48E"; 
		s_E585_C1_L				  :std_logic_vector(11 downto 0) := x"490"; 
		s_E586_C1_L				  :std_logic_vector(11 downto 0) := x"492"; 
		s_E587_C1_L				  :std_logic_vector(11 downto 0) := x"494"; 
		s_E588_C1_L				  :std_logic_vector(11 downto 0) := x"496"; 
		s_E589_C1_L				  :std_logic_vector(11 downto 0) := x"498"; 
		s_E590_C1_L				  :std_logic_vector(11 downto 0) := x"49A"; 
		s_E591_C1_L				  :std_logic_vector(11 downto 0) := x"49C"; 
		s_E592_C1_L				  :std_logic_vector(11 downto 0) := x"49E"; 
		s_E593_C1_L				  :std_logic_vector(11 downto 0) := x"4A0"; 
		s_E594_C1_L				  :std_logic_vector(11 downto 0) := x"4A2"; 
		s_E595_C1_L				  :std_logic_vector(11 downto 0) := x"4A4"; 
		s_E596_C1_L				  :std_logic_vector(11 downto 0) := x"4A6"; 
		s_E597_C1_L				  :std_logic_vector(11 downto 0) := x"4A8"; 
		s_E598_C1_L				  :std_logic_vector(11 downto 0) := x"4AA"; 
		s_E599_C1_L				  :std_logic_vector(11 downto 0) := x"4AC"; 
		s_E600_C1_L				  :std_logic_vector(11 downto 0) := x"4AE"; 
		s_E601_C1_L				  :std_logic_vector(11 downto 0) := x"4B0"; 
		s_E602_C1_L				  :std_logic_vector(11 downto 0) := x"4B2"; 
		s_E603_C1_L				  :std_logic_vector(11 downto 0) := x"4B4"; 
		s_E604_C1_L				  :std_logic_vector(11 downto 0) := x"4B6"; 
		s_E605_C1_L				  :std_logic_vector(11 downto 0) := x"4B8"; 
		s_E606_C1_L				  :std_logic_vector(11 downto 0) := x"4BA"; 
		s_E607_C1_L				  :std_logic_vector(11 downto 0) := x"4BC"; 
		s_E608_C1_L				  :std_logic_vector(11 downto 0) := x"4BE"; 
		s_E609_C1_L				  :std_logic_vector(11 downto 0) := x"4C0"; 
		s_E610_C1_L				  :std_logic_vector(11 downto 0) := x"4C2"; 
		s_E611_C1_L				  :std_logic_vector(11 downto 0) := x"4C4"; 
		s_E612_C1_L				  :std_logic_vector(11 downto 0) := x"4C6"; 
		s_E613_C1_L				  :std_logic_vector(11 downto 0) := x"4C8"; 
		s_E614_C1_L				  :std_logic_vector(11 downto 0) := x"4CA"; 
		s_E615_C1_L				  :std_logic_vector(11 downto 0) := x"4CC"; 
		s_E616_C1_L				  :std_logic_vector(11 downto 0) := x"4CE"; 
		s_E617_C1_L				  :std_logic_vector(11 downto 0) := x"4D0"; 
		s_E618_C1_L				  :std_logic_vector(11 downto 0) := x"4D2"; 
		s_E619_C1_L				  :std_logic_vector(11 downto 0) := x"4D4"; 
		s_E620_C1_L				  :std_logic_vector(11 downto 0) := x"4D6"; 
		s_E621_C1_L				  :std_logic_vector(11 downto 0) := x"4D8"; 
		s_E622_C1_L				  :std_logic_vector(11 downto 0) := x"4DA"; 
		s_E623_C1_L				  :std_logic_vector(11 downto 0) := x"4DC"; 
		s_E624_C1_L				  :std_logic_vector(11 downto 0) := x"4DE"; 
		s_E625_C1_L				  :std_logic_vector(11 downto 0) := x"4E0"; 
		s_E626_C1_L				  :std_logic_vector(11 downto 0) := x"4E2"; 
		s_E627_C1_L				  :std_logic_vector(11 downto 0) := x"4E4"; 
		s_E628_C1_L				  :std_logic_vector(11 downto 0) := x"4E6"; 
		s_E629_C1_L				  :std_logic_vector(11 downto 0) := x"4E8"; 
		s_E630_C1_L				  :std_logic_vector(11 downto 0) := x"4EA"; 
		s_E631_C1_L				  :std_logic_vector(11 downto 0) := x"4EC"; 
		s_E632_C1_L				  :std_logic_vector(11 downto 0) := x"4EE"; 
		s_E633_C1_L				  :std_logic_vector(11 downto 0) := x"4F0"; 
		s_E634_C1_L				  :std_logic_vector(11 downto 0) := x"4F2"; 
		s_E635_C1_L				  :std_logic_vector(11 downto 0) := x"4F4"; 
		s_E636_C1_L				  :std_logic_vector(11 downto 0) := x"4F6"; 
		s_E637_C1_L				  :std_logic_vector(11 downto 0) := x"4F8"; 
		s_E638_C1_L				  :std_logic_vector(11 downto 0) := x"4FA"; 
		s_E639_C1_L				  :std_logic_vector(11 downto 0) := x"4FC"; 
		s_E640_C1_L				  :std_logic_vector(11 downto 0) := x"4FE"; 
		s_E641_C1_L				  :std_logic_vector(11 downto 0) := x"500"; 
		s_E642_C1_L				  :std_logic_vector(11 downto 0) := x"502"; 
		s_E643_C1_L				  :std_logic_vector(11 downto 0) := x"504"; 
		s_E644_C1_L				  :std_logic_vector(11 downto 0) := x"506"; 
		s_E645_C1_L				  :std_logic_vector(11 downto 0) := x"508"; 
		s_E646_C1_L				  :std_logic_vector(11 downto 0) := x"50A"; 
		s_E647_C1_L				  :std_logic_vector(11 downto 0) := x"50C"; 
		s_E648_C1_L				  :std_logic_vector(11 downto 0) := x"50E"; 
		s_E649_C1_L				  :std_logic_vector(11 downto 0) := x"510"; 
		s_E650_C1_L				  :std_logic_vector(11 downto 0) := x"512"; 
		s_E651_C1_L				  :std_logic_vector(11 downto 0) := x"514"; 
		s_E652_C1_L				  :std_logic_vector(11 downto 0) := x"516"; 
		s_E653_C1_L				  :std_logic_vector(11 downto 0) := x"518"; 
		s_E654_C1_L				  :std_logic_vector(11 downto 0) := x"51A"; 
		s_E655_C1_L				  :std_logic_vector(11 downto 0) := x"51C"; 
		s_E656_C1_L				  :std_logic_vector(11 downto 0) := x"51E"; 
		s_E657_C1_L				  :std_logic_vector(11 downto 0) := x"520"; 
		s_E658_C1_L				  :std_logic_vector(11 downto 0) := x"522"; 
		s_E659_C1_L				  :std_logic_vector(11 downto 0) := x"524"; 
		s_E660_C1_L				  :std_logic_vector(11 downto 0) := x"526"; 
		s_E661_C1_L				  :std_logic_vector(11 downto 0) := x"528"; 
		s_E662_C1_L				  :std_logic_vector(11 downto 0) := x"52A"; 
		s_E663_C1_L				  :std_logic_vector(11 downto 0) := x"52C"; 
		s_E664_C1_L				  :std_logic_vector(11 downto 0) := x"52E"; 
		s_E665_C1_L				  :std_logic_vector(11 downto 0) := x"530"; 
		s_E666_C1_L				  :std_logic_vector(11 downto 0) := x"532"; 
		s_E667_C1_L				  :std_logic_vector(11 downto 0) := x"534"; 
		s_E668_C1_L				  :std_logic_vector(11 downto 0) := x"536"; 
		s_E669_C1_L				  :std_logic_vector(11 downto 0) := x"538"; 
		s_E670_C1_L				  :std_logic_vector(11 downto 0) := x"53A"; 
		s_E671_C1_L				  :std_logic_vector(11 downto 0) := x"53C"; 
		s_E672_C1_L				  :std_logic_vector(11 downto 0) := x"53E"; 
		s_E673_C1_L				  :std_logic_vector(11 downto 0) := x"540"; 
		s_E674_C1_L				  :std_logic_vector(11 downto 0) := x"542"; 
		s_E675_C1_L				  :std_logic_vector(11 downto 0) := x"544"; 
		s_E676_C1_L				  :std_logic_vector(11 downto 0) := x"546"; 
		s_E677_C1_L				  :std_logic_vector(11 downto 0) := x"548"; 
		s_E678_C1_L				  :std_logic_vector(11 downto 0) := x"54A"; 
		s_E679_C1_L				  :std_logic_vector(11 downto 0) := x"54C"; 
		s_E680_C1_L				  :std_logic_vector(11 downto 0) := x"54E"; 
		s_E681_C1_L				  :std_logic_vector(11 downto 0) := x"550"; 
		s_E682_C1_L				  :std_logic_vector(11 downto 0) := x"552"; 
		s_E683_C1_L				  :std_logic_vector(11 downto 0) := x"554"; 
		s_E684_C1_L				  :std_logic_vector(11 downto 0) := x"556"; 
		s_E685_C1_L				  :std_logic_vector(11 downto 0) := x"558"; 
		s_E686_C1_L				  :std_logic_vector(11 downto 0) := x"55A"; 
		s_E687_C1_L				  :std_logic_vector(11 downto 0) := x"55C"; 
		s_E688_C1_L				  :std_logic_vector(11 downto 0) := x"55E"; 
		s_E689_C1_L				  :std_logic_vector(11 downto 0) := x"560"; 
		s_E690_C1_L				  :std_logic_vector(11 downto 0) := x"562"; 
		s_E691_C1_L				  :std_logic_vector(11 downto 0) := x"564"; 
		s_E692_C1_L				  :std_logic_vector(11 downto 0) := x"566"; 
		s_E693_C1_L				  :std_logic_vector(11 downto 0) := x"568"; 
		s_E694_C1_L				  :std_logic_vector(11 downto 0) := x"56A"; 
		s_E695_C1_L				  :std_logic_vector(11 downto 0) := x"56C"; 
		s_E696_C1_L				  :std_logic_vector(11 downto 0) := x"56E"; 
		s_E697_C1_L				  :std_logic_vector(11 downto 0) := x"570"; 
		s_E698_C1_L				  :std_logic_vector(11 downto 0) := x"572"; 
		s_E699_C1_L				  :std_logic_vector(11 downto 0) := x"574"; 
		s_E700_C1_L				  :std_logic_vector(11 downto 0) := x"576"; 
		s_E701_C1_L				  :std_logic_vector(11 downto 0) := x"578"; 
		s_E702_C1_L				  :std_logic_vector(11 downto 0) := x"57A"; 
		s_E703_C1_L				  :std_logic_vector(11 downto 0) := x"57C"; 
		s_E704_C1_L				  :std_logic_vector(11 downto 0) := x"57E"; 
		s_E705_C1_L				  :std_logic_vector(11 downto 0) := x"580"; 
		s_E706_C1_L				  :std_logic_vector(11 downto 0) := x"582"; 
		s_E707_C1_L				  :std_logic_vector(11 downto 0) := x"584"; 
		s_E708_C1_L				  :std_logic_vector(11 downto 0) := x"586"; 
		s_E709_C1_L				  :std_logic_vector(11 downto 0) := x"588"; 
		s_E710_C1_L				  :std_logic_vector(11 downto 0) := x"58A"; 
		s_E711_C1_L				  :std_logic_vector(11 downto 0) := x"58C"; 
		s_E712_C1_L				  :std_logic_vector(11 downto 0) := x"58E"; 
		s_E713_C1_L				  :std_logic_vector(11 downto 0) := x"590"; 
		s_E714_C1_L				  :std_logic_vector(11 downto 0) := x"592"; 
		s_E715_C1_L				  :std_logic_vector(11 downto 0) := x"594"; 
		s_E716_C1_L				  :std_logic_vector(11 downto 0) := x"596"; 
		s_E717_C1_L				  :std_logic_vector(11 downto 0) := x"598"; 
		s_E718_C1_L				  :std_logic_vector(11 downto 0) := x"59A"; 
		s_E719_C1_L				  :std_logic_vector(11 downto 0) := x"59C"; 
		s_E720_C1_L				  :std_logic_vector(11 downto 0) := x"59E"; 
		s_E721_C1_L				  :std_logic_vector(11 downto 0) := x"5A0"; 
		s_E722_C1_L				  :std_logic_vector(11 downto 0) := x"5A2"; 
		s_E723_C1_L				  :std_logic_vector(11 downto 0) := x"5A4"; 
		s_E724_C1_L				  :std_logic_vector(11 downto 0) := x"5A6"; 
		s_E725_C1_L				  :std_logic_vector(11 downto 0) := x"5A8"; 
		s_E726_C1_L				  :std_logic_vector(11 downto 0) := x"5AA"; 
		s_E727_C1_L				  :std_logic_vector(11 downto 0) := x"5AC"; 
		s_E728_C1_L				  :std_logic_vector(11 downto 0) := x"5AE"; 
		s_E729_C1_L				  :std_logic_vector(11 downto 0) := x"5B0"; 
		s_E730_C1_L				  :std_logic_vector(11 downto 0) := x"5B2"; 
		s_E731_C1_L				  :std_logic_vector(11 downto 0) := x"5B4"; 
		s_E732_C1_L				  :std_logic_vector(11 downto 0) := x"5B6"; 
		s_E733_C1_L				  :std_logic_vector(11 downto 0) := x"5B8"; 
		s_E734_C1_L				  :std_logic_vector(11 downto 0) := x"5BA"; 
		s_E735_C1_L				  :std_logic_vector(11 downto 0) := x"5BC"; 
		s_E736_C1_L				  :std_logic_vector(11 downto 0) := x"5BE"; 
		s_E737_C1_L				  :std_logic_vector(11 downto 0) := x"5C0"; 
		s_E738_C1_L				  :std_logic_vector(11 downto 0) := x"5C2"; 
		s_E739_C1_L				  :std_logic_vector(11 downto 0) := x"5C4"; 
		s_E740_C1_L				  :std_logic_vector(11 downto 0) := x"5C6"; 
		s_E741_C1_L				  :std_logic_vector(11 downto 0) := x"5C8"; 
		s_E742_C1_L				  :std_logic_vector(11 downto 0) := x"5CA"; 
		s_E743_C1_L				  :std_logic_vector(11 downto 0) := x"5CC"; 
		s_E744_C1_L				  :std_logic_vector(11 downto 0) := x"5CE"; 
		s_E745_C1_L				  :std_logic_vector(11 downto 0) := x"5D0"; 
		s_E746_C1_L				  :std_logic_vector(11 downto 0) := x"5D2"; 
		s_E747_C1_L				  :std_logic_vector(11 downto 0) := x"5D4"; 
		s_E748_C1_L				  :std_logic_vector(11 downto 0) := x"5D6"; 
		s_E749_C1_L				  :std_logic_vector(11 downto 0) := x"5D8"; 
		s_E750_C1_L				  :std_logic_vector(11 downto 0) := x"5DA"; 
		s_E751_C1_L				  :std_logic_vector(11 downto 0) := x"5DC"; 
		s_E752_C1_L				  :std_logic_vector(11 downto 0) := x"5DE"; 
		s_E753_C1_L				  :std_logic_vector(11 downto 0) := x"5E0"; 
		s_E754_C1_L				  :std_logic_vector(11 downto 0) := x"5E2"; 
		s_E755_C1_L				  :std_logic_vector(11 downto 0) := x"5E4"; 
		s_E756_C1_L				  :std_logic_vector(11 downto 0) := x"5E6"; 
		s_E757_C1_L				  :std_logic_vector(11 downto 0) := x"5E8"; 
		s_E758_C1_L				  :std_logic_vector(11 downto 0) := x"5EA"; 
		s_E759_C1_L				  :std_logic_vector(11 downto 0) := x"5EC"; 
		s_E760_C1_L				  :std_logic_vector(11 downto 0) := x"5EE"; 
		s_E761_C1_L				  :std_logic_vector(11 downto 0) := x"5F0"; 
		s_E762_C1_L				  :std_logic_vector(11 downto 0) := x"5F2"; 
		s_E763_C1_L				  :std_logic_vector(11 downto 0) := x"5F4"; 
		s_E764_C1_L				  :std_logic_vector(11 downto 0) := x"5F6"; 
		s_E765_C1_L				  :std_logic_vector(11 downto 0) := x"5F8"; 
		s_E766_C1_L				  :std_logic_vector(11 downto 0) := x"5FA"; 
		s_E767_C1_L				  :std_logic_vector(11 downto 0) := x"5FC"; 
		s_E768_C1_L				  :std_logic_vector(11 downto 0) := x"5FE"; 
		s_E769_C1_L				  :std_logic_vector(11 downto 0) := x"600"; 
		s_E770_C1_L				  :std_logic_vector(11 downto 0) := x"602"; 
		s_E771_C1_L				  :std_logic_vector(11 downto 0) := x"604"; 
		s_E772_C1_L				  :std_logic_vector(11 downto 0) := x"606"; 
		s_E773_C1_L				  :std_logic_vector(11 downto 0) := x"608"; 
		s_E774_C1_L				  :std_logic_vector(11 downto 0) := x"60A"; 
		s_E775_C1_L				  :std_logic_vector(11 downto 0) := x"60C"; 
		s_E776_C1_L				  :std_logic_vector(11 downto 0) := x"60E"; 
		s_E777_C1_L				  :std_logic_vector(11 downto 0) := x"610"; 
		s_E778_C1_L				  :std_logic_vector(11 downto 0) := x"612"; 
		s_E779_C1_L				  :std_logic_vector(11 downto 0) := x"614"; 
		s_E780_C1_L				  :std_logic_vector(11 downto 0) := x"616"; 
		s_E781_C1_L				  :std_logic_vector(11 downto 0) := x"618"; 
		s_E782_C1_L				  :std_logic_vector(11 downto 0) := x"61A"; 
		s_E783_C1_L				  :std_logic_vector(11 downto 0) := x"61C"; 
		s_E784_C1_L				  :std_logic_vector(11 downto 0) := x"61E"; 
		s_E785_C1_L				  :std_logic_vector(11 downto 0) := x"620"; 
		s_E786_C1_L				  :std_logic_vector(11 downto 0) := x"622"; 
		s_E787_C1_L				  :std_logic_vector(11 downto 0) := x"624"; 
		s_E788_C1_L				  :std_logic_vector(11 downto 0) := x"626"; 
		s_E789_C1_L				  :std_logic_vector(11 downto 0) := x"628"; 
		s_E790_C1_L				  :std_logic_vector(11 downto 0) := x"62A"; 
		s_E791_C1_L				  :std_logic_vector(11 downto 0) := x"62C"; 
		s_E792_C1_L				  :std_logic_vector(11 downto 0) := x"62E"; 
		s_E793_C1_L				  :std_logic_vector(11 downto 0) := x"630"; 
		s_E794_C1_L				  :std_logic_vector(11 downto 0) := x"632"; 
		s_E795_C1_L				  :std_logic_vector(11 downto 0) := x"634"; 
		s_E796_C1_L				  :std_logic_vector(11 downto 0) := x"636"; 
		s_E797_C1_L				  :std_logic_vector(11 downto 0) := x"638"; 
		s_E798_C1_L				  :std_logic_vector(11 downto 0) := x"63A"; 
		s_E799_C1_L				  :std_logic_vector(11 downto 0) := x"63C"; 
		s_E800_C1_L				  :std_logic_vector(11 downto 0) := x"63E"; 
		s_E801_C1_L				  :std_logic_vector(11 downto 0) := x"640"; 
		s_E802_C1_L				  :std_logic_vector(11 downto 0) := x"642"; 
		s_E803_C1_L				  :std_logic_vector(11 downto 0) := x"644"; 
		s_E804_C1_L				  :std_logic_vector(11 downto 0) := x"646"; 
		s_E805_C1_L				  :std_logic_vector(11 downto 0) := x"648"; 
		s_E806_C1_L				  :std_logic_vector(11 downto 0) := x"64A"; 
		s_E807_C1_L				  :std_logic_vector(11 downto 0) := x"64C"; 
		s_E808_C1_L				  :std_logic_vector(11 downto 0) := x"64E"; 
		s_E809_C1_L				  :std_logic_vector(11 downto 0) := x"650"; 
		s_E810_C1_L				  :std_logic_vector(11 downto 0) := x"652"; 
		s_E811_C1_L				  :std_logic_vector(11 downto 0) := x"654"; 
		s_E812_C1_L				  :std_logic_vector(11 downto 0) := x"656"; 
		s_E813_C1_L				  :std_logic_vector(11 downto 0) := x"658"; 
		s_E814_C1_L				  :std_logic_vector(11 downto 0) := x"65A"; 
		s_E815_C1_L				  :std_logic_vector(11 downto 0) := x"65C"; 
		s_E816_C1_L				  :std_logic_vector(11 downto 0) := x"65E"; 
		s_E817_C1_L				  :std_logic_vector(11 downto 0) := x"660"; 
		s_E818_C1_L				  :std_logic_vector(11 downto 0) := x"662"; 
		s_E819_C1_L				  :std_logic_vector(11 downto 0) := x"664"; 
		s_E820_C1_L				  :std_logic_vector(11 downto 0) := x"666"; 
		s_E821_C1_L				  :std_logic_vector(11 downto 0) := x"668"; 
		s_E822_C1_L				  :std_logic_vector(11 downto 0) := x"66A"; 
		s_E823_C1_L				  :std_logic_vector(11 downto 0) := x"66C"; 
		s_E824_C1_L				  :std_logic_vector(11 downto 0) := x"66E"; 
		s_E825_C1_L				  :std_logic_vector(11 downto 0) := x"670"; 
		s_E826_C1_L				  :std_logic_vector(11 downto 0) := x"672"; 
		s_E827_C1_L				  :std_logic_vector(11 downto 0) := x"674"; 
		s_E828_C1_L				  :std_logic_vector(11 downto 0) := x"676"; 
		s_E829_C1_L				  :std_logic_vector(11 downto 0) := x"678"; 
		s_E830_C1_L				  :std_logic_vector(11 downto 0) := x"67A"; 
		s_E831_C1_L				  :std_logic_vector(11 downto 0) := x"67C"; 
		s_E832_C1_L				  :std_logic_vector(11 downto 0) := x"67E"; 
		s_E833_C1_L				  :std_logic_vector(11 downto 0) := x"680"; 
		s_E834_C1_L				  :std_logic_vector(11 downto 0) := x"682"; 
		s_E835_C1_L				  :std_logic_vector(11 downto 0) := x"684"; 
		s_E836_C1_L				  :std_logic_vector(11 downto 0) := x"686"; 
		s_E837_C1_L				  :std_logic_vector(11 downto 0) := x"688"; 
		s_E838_C1_L				  :std_logic_vector(11 downto 0) := x"68A"; 
		s_E839_C1_L				  :std_logic_vector(11 downto 0) := x"68C"; 
		s_E840_C1_L				  :std_logic_vector(11 downto 0) := x"68E"; 
		s_E841_C1_L				  :std_logic_vector(11 downto 0) := x"690"; 
		s_E842_C1_L				  :std_logic_vector(11 downto 0) := x"692"; 
		s_E843_C1_L				  :std_logic_vector(11 downto 0) := x"694"; 
		s_E844_C1_L				  :std_logic_vector(11 downto 0) := x"696"; 
		s_E845_C1_L				  :std_logic_vector(11 downto 0) := x"698"; 
		s_E846_C1_L				  :std_logic_vector(11 downto 0) := x"69A"; 
		s_E847_C1_L				  :std_logic_vector(11 downto 0) := x"69C"; 
		s_E848_C1_L				  :std_logic_vector(11 downto 0) := x"69E"; 
		s_E849_C1_L				  :std_logic_vector(11 downto 0) := x"6A0"; 
		s_E850_C1_L				  :std_logic_vector(11 downto 0) := x"6A2"; 
		s_E851_C1_L				  :std_logic_vector(11 downto 0) := x"6A4"; 
		s_E852_C1_L				  :std_logic_vector(11 downto 0) := x"6A6"; 
		s_E853_C1_L				  :std_logic_vector(11 downto 0) := x"6A8"; 
		s_E854_C1_L				  :std_logic_vector(11 downto 0) := x"6AA"; 
		s_E855_C1_L				  :std_logic_vector(11 downto 0) := x"6AC"; 
		s_E856_C1_L				  :std_logic_vector(11 downto 0) := x"6AE"; 
		s_E857_C1_L				  :std_logic_vector(11 downto 0) := x"6B0"; 
		s_E858_C1_L				  :std_logic_vector(11 downto 0) := x"6B2"; 
		s_E859_C1_L				  :std_logic_vector(11 downto 0) := x"6B4"; 
		s_E860_C1_L				  :std_logic_vector(11 downto 0) := x"6B6"; 
		s_E861_C1_L				  :std_logic_vector(11 downto 0) := x"6B8"; 
		s_E862_C1_L				  :std_logic_vector(11 downto 0) := x"6BA"; 
		s_E863_C1_L				  :std_logic_vector(11 downto 0) := x"6BC"; 
		s_E864_C1_L				  :std_logic_vector(11 downto 0) := x"6BE"; 
		s_E865_C1_L				  :std_logic_vector(11 downto 0) := x"6C0"; 
		s_E866_C1_L				  :std_logic_vector(11 downto 0) := x"6C2"; 
		s_E867_C1_L				  :std_logic_vector(11 downto 0) := x"6C4"; 
		s_E868_C1_L				  :std_logic_vector(11 downto 0) := x"6C6"; 
		s_E869_C1_L				  :std_logic_vector(11 downto 0) := x"6C8"; 
		s_E870_C1_L				  :std_logic_vector(11 downto 0) := x"6CA"; 
		s_E871_C1_L				  :std_logic_vector(11 downto 0) := x"6CC"; 
		s_E872_C1_L				  :std_logic_vector(11 downto 0) := x"6CE"; 
		s_E873_C1_L				  :std_logic_vector(11 downto 0) := x"6D0"; 
		s_E874_C1_L				  :std_logic_vector(11 downto 0) := x"6D2"; 
		s_E875_C1_L				  :std_logic_vector(11 downto 0) := x"6D4"; 
		s_E876_C1_L				  :std_logic_vector(11 downto 0) := x"6D6"; 
		s_E877_C1_L				  :std_logic_vector(11 downto 0) := x"6D8"; 
		s_E878_C1_L				  :std_logic_vector(11 downto 0) := x"6DA"; 
		s_E879_C1_L				  :std_logic_vector(11 downto 0) := x"6DC"; 
		s_E880_C1_L				  :std_logic_vector(11 downto 0) := x"6DE"; 
		s_E881_C1_L				  :std_logic_vector(11 downto 0) := x"6E0"; 
		s_E882_C1_L				  :std_logic_vector(11 downto 0) := x"6E2"; 
		s_E883_C1_L				  :std_logic_vector(11 downto 0) := x"6E4"; 
		s_E884_C1_L				  :std_logic_vector(11 downto 0) := x"6E6"; 
		s_E885_C1_L				  :std_logic_vector(11 downto 0) := x"6E8"; 
		s_E886_C1_L				  :std_logic_vector(11 downto 0) := x"6EA"; 
		s_E887_C1_L				  :std_logic_vector(11 downto 0) := x"6EC"; 
		s_E888_C1_L				  :std_logic_vector(11 downto 0) := x"6EE"; 
		s_E889_C1_L				  :std_logic_vector(11 downto 0) := x"6F0"; 
		s_E890_C1_L				  :std_logic_vector(11 downto 0) := x"6F2"; 
		s_E891_C1_L				  :std_logic_vector(11 downto 0) := x"6F4"; 
		s_E892_C1_L				  :std_logic_vector(11 downto 0) := x"6F6"; 
		s_E893_C1_L				  :std_logic_vector(11 downto 0) := x"6F8"; 
		s_E894_C1_L				  :std_logic_vector(11 downto 0) := x"6FA"; 
		s_E895_C1_L				  :std_logic_vector(11 downto 0) := x"6FC"; 
		s_E896_C1_L				  :std_logic_vector(11 downto 0) := x"6FE"; 
		s_E897_C1_L				  :std_logic_vector(11 downto 0) := x"700"; 
		s_E898_C1_L				  :std_logic_vector(11 downto 0) := x"702"; 
		s_E899_C1_L				  :std_logic_vector(11 downto 0) := x"704"; 
		s_E900_C1_L				  :std_logic_vector(11 downto 0) := x"706"; 
		s_E901_C1_L				  :std_logic_vector(11 downto 0) := x"708"; 
		s_E902_C1_L				  :std_logic_vector(11 downto 0) := x"70A"; 
		s_E903_C1_L				  :std_logic_vector(11 downto 0) := x"70C"; 
		s_E904_C1_L				  :std_logic_vector(11 downto 0) := x"70E"; 
		s_E905_C1_L				  :std_logic_vector(11 downto 0) := x"710"; 
		s_E906_C1_L				  :std_logic_vector(11 downto 0) := x"712"; 
		s_E907_C1_L				  :std_logic_vector(11 downto 0) := x"714"; 
		s_E908_C1_L				  :std_logic_vector(11 downto 0) := x"716"; 
		s_E909_C1_L				  :std_logic_vector(11 downto 0) := x"718"; 
		s_E910_C1_L				  :std_logic_vector(11 downto 0) := x"71A"; 
		s_E911_C1_L				  :std_logic_vector(11 downto 0) := x"71C"; 
		s_E912_C1_L				  :std_logic_vector(11 downto 0) := x"71E"; 
		s_E913_C1_L				  :std_logic_vector(11 downto 0) := x"720"; 
		s_E914_C1_L				  :std_logic_vector(11 downto 0) := x"722"; 
		s_E915_C1_L				  :std_logic_vector(11 downto 0) := x"724"; 
		s_E916_C1_L				  :std_logic_vector(11 downto 0) := x"726"; 
		s_E917_C1_L				  :std_logic_vector(11 downto 0) := x"728"; 
		s_E918_C1_L				  :std_logic_vector(11 downto 0) := x"72A"; 
		s_E919_C1_L				  :std_logic_vector(11 downto 0) := x"72C"; 
		s_E920_C1_L				  :std_logic_vector(11 downto 0) := x"72E"; 
		s_E921_C1_L				  :std_logic_vector(11 downto 0) := x"730"; 
		s_E922_C1_L				  :std_logic_vector(11 downto 0) := x"732"; 
		s_E923_C1_L				  :std_logic_vector(11 downto 0) := x"734"; 
		s_E924_C1_L				  :std_logic_vector(11 downto 0) := x"736"; 
		s_E925_C1_L				  :std_logic_vector(11 downto 0) := x"738"; 
		s_E926_C1_L				  :std_logic_vector(11 downto 0) := x"73A"; 
		s_E927_C1_L				  :std_logic_vector(11 downto 0) := x"73C"; 
		s_E928_C1_L				  :std_logic_vector(11 downto 0) := x"73E"; 
		s_E929_C1_L				  :std_logic_vector(11 downto 0) := x"740"; 
		s_E930_C1_L				  :std_logic_vector(11 downto 0) := x"742"; 
		s_E931_C1_L				  :std_logic_vector(11 downto 0) := x"744"; 
		s_E932_C1_L				  :std_logic_vector(11 downto 0) := x"746"; 
		s_E933_C1_L				  :std_logic_vector(11 downto 0) := x"748"; 
		s_E934_C1_L				  :std_logic_vector(11 downto 0) := x"74A"; 
		s_E935_C1_L				  :std_logic_vector(11 downto 0) := x"74C"; 
		s_E936_C1_L				  :std_logic_vector(11 downto 0) := x"74E"; 
		s_E937_C1_L				  :std_logic_vector(11 downto 0) := x"750"; 
		s_E938_C1_L				  :std_logic_vector(11 downto 0) := x"752"; 
		s_E939_C1_L				  :std_logic_vector(11 downto 0) := x"754"; 
		s_E940_C1_L				  :std_logic_vector(11 downto 0) := x"756"; 
		s_E941_C1_L				  :std_logic_vector(11 downto 0) := x"758"; 
		s_E942_C1_L				  :std_logic_vector(11 downto 0) := x"75A"; 
		s_E943_C1_L				  :std_logic_vector(11 downto 0) := x"75C"; 
		s_E944_C1_L				  :std_logic_vector(11 downto 0) := x"75E"; 
		s_E945_C1_L				  :std_logic_vector(11 downto 0) := x"760"; 
		s_E946_C1_L				  :std_logic_vector(11 downto 0) := x"762"; 
		s_E947_C1_L				  :std_logic_vector(11 downto 0) := x"764"; 
		s_E948_C1_L				  :std_logic_vector(11 downto 0) := x"766"; 
		s_E949_C1_L				  :std_logic_vector(11 downto 0) := x"768"; 
		s_E950_C1_L				  :std_logic_vector(11 downto 0) := x"76A"; 
		s_E951_C1_L				  :std_logic_vector(11 downto 0) := x"76C"; 
		s_E952_C1_L				  :std_logic_vector(11 downto 0) := x"76E"; 
		s_E953_C1_L				  :std_logic_vector(11 downto 0) := x"770"; 
		s_E954_C1_L				  :std_logic_vector(11 downto 0) := x"772"; 
		s_E955_C1_L				  :std_logic_vector(11 downto 0) := x"774"; 
		s_E956_C1_L				  :std_logic_vector(11 downto 0) := x"776"; 
		s_E957_C1_L				  :std_logic_vector(11 downto 0) := x"778"; 
		s_E958_C1_L				  :std_logic_vector(11 downto 0) := x"77A"; 
		s_E959_C1_L				  :std_logic_vector(11 downto 0) := x"77C"; 
		s_E960_C1_L				  :std_logic_vector(11 downto 0) := x"77E"; 
		s_E961_C1_L				  :std_logic_vector(11 downto 0) := x"780"; 
		s_E962_C1_L				  :std_logic_vector(11 downto 0) := x"782"; 
		s_E963_C1_L				  :std_logic_vector(11 downto 0) := x"784"; 
		s_E964_C1_L				  :std_logic_vector(11 downto 0) := x"786"; 
		s_E965_C1_L				  :std_logic_vector(11 downto 0) := x"788"; 
		s_E966_C1_L				  :std_logic_vector(11 downto 0) := x"78A"; 
		s_E967_C1_L				  :std_logic_vector(11 downto 0) := x"78C"; 
		s_E968_C1_L				  :std_logic_vector(11 downto 0) := x"78E"; 
		s_E969_C1_L				  :std_logic_vector(11 downto 0) := x"790"; 
		s_E970_C1_L				  :std_logic_vector(11 downto 0) := x"792"; 
		s_E971_C1_L				  :std_logic_vector(11 downto 0) := x"794"; 
		s_E972_C1_L				  :std_logic_vector(11 downto 0) := x"796"; 
		s_E973_C1_L				  :std_logic_vector(11 downto 0) := x"798"; 
		s_E974_C1_L				  :std_logic_vector(11 downto 0) := x"79A"; 
		s_E975_C1_L				  :std_logic_vector(11 downto 0) := x"79C"; 
		s_E976_C1_L				  :std_logic_vector(11 downto 0) := x"79E"; 
		s_E977_C1_L				  :std_logic_vector(11 downto 0) := x"7A0"; 
		s_E978_C1_L				  :std_logic_vector(11 downto 0) := x"7A2"; 
		s_E979_C1_L				  :std_logic_vector(11 downto 0) := x"7A4"; 
		s_E980_C1_L				  :std_logic_vector(11 downto 0) := x"7A6"; 
		s_E981_C1_L				  :std_logic_vector(11 downto 0) := x"7A8"; 
		s_E982_C1_L				  :std_logic_vector(11 downto 0) := x"7AA"; 
		s_E983_C1_L				  :std_logic_vector(11 downto 0) := x"7AC"; 
		s_E984_C1_L				  :std_logic_vector(11 downto 0) := x"7AE"; 
		s_E985_C1_L				  :std_logic_vector(11 downto 0) := x"7B0"; 
		s_E986_C1_L				  :std_logic_vector(11 downto 0) := x"7B2"; 
		s_E987_C1_L				  :std_logic_vector(11 downto 0) := x"7B4"; 
		s_E988_C1_L				  :std_logic_vector(11 downto 0) := x"7B6"; 
		s_E989_C1_L				  :std_logic_vector(11 downto 0) := x"7B8"; 
		s_E990_C1_L				  :std_logic_vector(11 downto 0) := x"7BA"; 
		s_E991_C1_L				  :std_logic_vector(11 downto 0) := x"7BC"; 
		s_E992_C1_L				  :std_logic_vector(11 downto 0) := x"7BE"; 
		s_E993_C1_L				  :std_logic_vector(11 downto 0) := x"7C0"; 
		s_E994_C1_L				  :std_logic_vector(11 downto 0) := x"7C2"; 
		s_E995_C1_L				  :std_logic_vector(11 downto 0) := x"7C4"; 
		s_E996_C1_L				  :std_logic_vector(11 downto 0) := x"7C6"; 
		s_E997_C1_L				  :std_logic_vector(11 downto 0) := x"7C8"; 
		s_E998_C1_L				  :std_logic_vector(11 downto 0) := x"7CA"; 
		s_E999_C1_L				  :std_logic_vector(11 downto 0) := x"7CC"; 
		s_E1000_C1_L			  :std_logic_vector(11 downto 0) := x"7CE"; 
		s_E1001_C1_L			  :std_logic_vector(11 downto 0) := x"7D0"; 
		s_E1002_C1_L			  :std_logic_vector(11 downto 0) := x"7D2"; 
		s_E1003_C1_L			  :std_logic_vector(11 downto 0) := x"7D4"; 
		s_E1004_C1_L			  :std_logic_vector(11 downto 0) := x"7D6"; 
		s_E1005_C1_L			  :std_logic_vector(11 downto 0) := x"7D8"; 
		s_E1006_C1_L			  :std_logic_vector(11 downto 0) := x"7DA"; 
		s_E1007_C1_L			  :std_logic_vector(11 downto 0) := x"7DC"; 
		s_E1008_C1_L			  :std_logic_vector(11 downto 0) := x"7DE"; 
		s_E1009_C1_L			  :std_logic_vector(11 downto 0) := x"7E0"; 
		s_E1010_C1_L			  :std_logic_vector(11 downto 0) := x"7E2"; 
		s_E1011_C1_L			  :std_logic_vector(11 downto 0) := x"7E4"; 
		s_E1012_C1_L			  :std_logic_vector(11 downto 0) := x"7E6"; 
		s_E1013_C1_L			  :std_logic_vector(11 downto 0) := x"7E8"; 
		s_E1014_C1_L			  :std_logic_vector(11 downto 0) := x"7EA"; 
		s_E1015_C1_L			  :std_logic_vector(11 downto 0) := x"7EC"; 
		s_E1016_C1_L			  :std_logic_vector(11 downto 0) := x"7EE"; 
		s_E1017_C1_L			  :std_logic_vector(11 downto 0) := x"7F0"; 
		s_E1018_C1_L			  :std_logic_vector(11 downto 0) := x"7F2"; 
		s_E1019_C1_L			  :std_logic_vector(11 downto 0) := x"7F4"; 
		s_E1020_C1_L			  :std_logic_vector(11 downto 0) := x"7F6"; 
		s_E1021_C1_L			  :std_logic_vector(11 downto 0) := x"7F8"; 
		s_E1022_C1_L			  :std_logic_vector(11 downto 0) := x"7FA"; 
		s_E1023_C1_L			  :std_logic_vector(11 downto 0) := x"7FC"; 
		s_E1024_C1_L			  :std_logic_vector(11 downto 0) := x"7FE"; 
                                                                    
		s_E1_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"7FF";
		s_E1_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"801";
		s_E2_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"803";
		s_E3_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"805";
		s_E4_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"807";
		s_E5_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"809";
		s_E6_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"80B";
		s_E7_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"80D";
		s_E8_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"80F";
		s_E9_C1_H_Pos        	  :std_logic_vector(11 downto 0) := x"811";
		s_E10_C1_H_Pos       	  :std_logic_vector(11 downto 0) := x"813";
		s_E11_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"815";
		s_E12_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"817";
		s_E13_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"819";
		s_E14_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"81B";
		s_E15_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"81D";
		s_E16_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"81F";
		s_E17_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"821";
		s_E18_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"823";
		s_E19_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"825";
		s_E20_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"827";
		s_E21_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"829";
		s_E22_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"82B";
		s_E23_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"82D";
		s_E24_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"82F";
		s_E25_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"831";
		s_E26_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"833";
		s_E27_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"835";
		s_E28_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"837";
		s_E29_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"839";
		s_E30_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"83B";
		s_E31_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"83D";
		s_E32_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"83F";
		s_E33_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"841";
		s_E34_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"843";
		s_E35_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"845";
		s_E36_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"847";
		s_E37_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"849";
		s_E38_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"84B";
		s_E39_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"84D";
		s_E40_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"84F";
		s_E41_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"851";
		s_E42_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"853";
		s_E43_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"855";
		s_E44_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"857";
		s_E45_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"859";
		s_E46_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"85B";
		s_E47_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"85D";
		s_E48_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"85F";
		s_E49_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"861";
		s_E50_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"863";
		s_E51_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"865";
		s_E52_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"867";
		s_E53_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"869";
		s_E54_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"86B";
		s_E55_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"86D";
		s_E56_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"86F";
		s_E57_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"871";
		s_E58_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"873";
		s_E59_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"875";
		s_E60_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"877";
		s_E61_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"879";
		s_E62_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"87B";
		s_E63_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"87D";
		s_E64_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"87F";
		s_E65_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"881";
		s_E66_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"883";
		s_E67_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"885";
		s_E68_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"887";
		s_E69_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"889";
		s_E70_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"88B";
		s_E71_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"88D";
		s_E72_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"88F";
		s_E73_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"891";
		s_E74_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"893";
		s_E75_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"895";
		s_E76_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"897";
		s_E77_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"899";
		s_E78_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"89B";
		s_E79_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"89D";
		s_E80_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"89F";
		s_E81_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8A1";
		s_E82_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8A3";
		s_E83_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8A5";
		s_E84_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8A7";
		s_E85_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8A9";
		s_E86_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8AB";
		s_E87_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8AD";
		s_E88_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8AF";
		s_E89_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8B1";
		s_E90_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8B3";
		s_E91_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8B5";
		s_E92_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8B7";
		s_E93_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8B9";
		s_E94_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8BB";
		s_E95_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8BD";
		s_E96_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8BF";
		s_E97_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8C1";
		s_E98_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8C3";
		s_E99_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8C5";
		s_E100_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8C7";
		s_E101_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8C9";
		s_E102_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8CB";
		s_E103_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8CD";
		s_E104_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8CF";
		s_E105_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8D1";
		s_E106_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8D3";
		s_E107_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8D5";
		s_E108_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8D7";
		s_E109_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8D9";
		s_E110_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8DB";
		s_E111_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8DD";
		s_E112_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8DF";
		s_E113_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8E1";
		s_E114_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8E3";
		s_E115_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8E5";
		s_E116_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8E7";
		s_E117_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8E9";
		s_E118_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8EB";
		s_E119_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8ED";
		s_E120_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8EF";
		s_E121_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8F1";
		s_E122_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8F3";
		s_E123_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8F5";
		s_E124_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8F7";
		s_E125_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8F9";
		s_E126_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8FB";
		s_E127_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8FD";
		s_E128_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"8FF";
		s_E129_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"901";
		s_E130_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"903";
		s_E131_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"905";
		s_E132_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"907";
		s_E133_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"909";
		s_E134_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"90B";
		s_E135_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"90D";
		s_E136_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"90F";
		s_E137_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"911";
		s_E138_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"913";
		s_E139_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"915";
		s_E140_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"917";
		s_E141_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"919";
		s_E142_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"91B";
		s_E143_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"91D";
		s_E144_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"91F";
		s_E145_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"921";
		s_E146_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"923";
		s_E147_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"925";
		s_E148_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"927";
		s_E149_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"929";
		s_E150_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"92B";
		s_E151_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"92D";
		s_E152_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"92F";
		s_E153_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"931";
		s_E154_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"933";
		s_E155_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"935";
		s_E156_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"937";
		s_E157_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"939";
		s_E158_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"93B";
		s_E159_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"93D";
		s_E160_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"93F";
		s_E161_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"941";
		s_E162_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"943";
		s_E163_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"945";
		s_E164_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"947";
		s_E165_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"949";
		s_E166_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"94B";
		s_E167_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"94D";
		s_E168_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"94F";
		s_E169_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"951";
		s_E170_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"953";
		s_E171_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"955";
		s_E172_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"957";
		s_E173_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"959";
		s_E174_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"95B";
		s_E175_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"95D";
		s_E176_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"95F";
		s_E177_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"961";
		s_E178_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"963";
		s_E179_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"965";
		s_E180_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"967";
		s_E181_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"969";
		s_E182_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"96B";
		s_E183_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"96D";
		s_E184_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"96F";
		s_E185_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"971";
		s_E186_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"973";
		s_E187_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"975";
		s_E188_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"977";
		s_E189_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"979";
		s_E190_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"97B";
		s_E191_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"97D";
		s_E192_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"97F";
		s_E193_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"981";
		s_E194_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"983";
		s_E195_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"985";
		s_E196_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"987";
		s_E197_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"989";
		s_E198_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"98B";
		s_E199_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"98D";
		s_E200_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"98F";
		s_E201_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"991";
		s_E202_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"993";
		s_E203_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"995";
		s_E204_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"997";
		s_E205_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"999";
		s_E206_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"99B";
		s_E207_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"99D";
		s_E208_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"99F";
		s_E209_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9A1";
		s_E210_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9A3";
		s_E211_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9A5";
		s_E212_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9A7";
		s_E213_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9A9";
		s_E214_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9AB";
		s_E215_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9AD";
		s_E216_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9AF";
		s_E217_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9B1";
		s_E218_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9B3";
		s_E219_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9B5";
		s_E220_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9B7";
		s_E221_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9B9";
		s_E222_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9BB";
		s_E223_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9BD";
		s_E224_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9BF";
		s_E225_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9C1";
		s_E226_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9C3";
		s_E227_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9C5";
		s_E228_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9C7";
		s_E229_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9C9";
		s_E230_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9CB";
		s_E231_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9CD";
		s_E232_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9CF";
		s_E233_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9D1";
		s_E234_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9D3";
		s_E235_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9D5";
		s_E236_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9D7";
		s_E237_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9D9";
		s_E238_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9DB";
		s_E239_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9DD";
		s_E240_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9DF";
		s_E241_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9E1";
		s_E242_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9E3";
		s_E243_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9E5";
		s_E244_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9E7";
		s_E245_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9E9";
		s_E246_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9EB";
		s_E247_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9ED";
		s_E248_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9EF";
		s_E249_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9F1";
		s_E250_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9F3";
		s_E251_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9F5";
		s_E252_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9F7";
		s_E253_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9F9";
		s_E254_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9FB";
		s_E255_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9FD";
		s_E256_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"9FF";
		s_E257_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A01";
		s_E258_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A03";
		s_E259_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A05";
		s_E260_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A07";
		s_E261_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A09";
		s_E262_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A0B";
		s_E263_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A0D";
		s_E264_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A0F";
		s_E265_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A11";
		s_E266_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A13";
		s_E267_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A15";
		s_E268_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A17";
		s_E269_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A19";
		s_E270_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A1B";
		s_E271_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A1D";
		s_E272_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A1F";
		s_E273_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A21";
		s_E274_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A23";
		s_E275_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A25";
		s_E276_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A27";
		s_E277_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A29";
		s_E278_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A2B";
		s_E279_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A2D";
		s_E280_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A2F";
		s_E281_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A31";
		s_E282_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A33";
		s_E283_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A35";
		s_E284_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A37";
		s_E285_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A39";
		s_E286_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A3B";
		s_E287_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A3D";
		s_E288_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A3F";
		s_E289_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A41";
		s_E290_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A43";
		s_E291_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A45";
		s_E292_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A47";
		s_E293_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A49";
		s_E294_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A4B";
		s_E295_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A4D";
		s_E296_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A4F";
		s_E297_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A51";
		s_E298_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A53";
		s_E299_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A55";
		s_E300_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A57";
		s_E301_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A59";
		s_E302_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A5B";
		s_E303_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A5D";
		s_E304_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A5F";
		s_E305_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A61";
		s_E306_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A63";
		s_E307_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A65";
		s_E308_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A67";
		s_E309_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A69";
		s_E310_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A6B";
		s_E311_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A6D";
		s_E312_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A6F";
		s_E313_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A71";
		s_E314_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A73";
		s_E315_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A75";
		s_E316_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A77";
		s_E317_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A79";
		s_E318_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A7B";
		s_E319_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A7D";
		s_E320_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A7F";
		s_E321_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A81";
		s_E322_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A83";
		s_E323_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A85";
		s_E324_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A87";
		s_E325_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A89";
		s_E326_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A8B";
		s_E327_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A8D";
		s_E328_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A8F";
		s_E329_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A91";
		s_E330_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A93";
		s_E331_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A95";
		s_E332_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A97";
		s_E333_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A99";
		s_E334_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A9B";
		s_E335_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A9D";
		s_E336_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"A9F";
		s_E337_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AA1";
		s_E338_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AA3";
		s_E339_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AA5";
		s_E340_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AA7";
		s_E341_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AA9";
		s_E342_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AAB";
		s_E343_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AAD";
		s_E344_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AAF";
		s_E345_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AB1";
		s_E346_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AB3";
		s_E347_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AB5";
		s_E348_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AB7";
		s_E349_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AB9";
		s_E350_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ABB";
		s_E351_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ABD";
		s_E352_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ABF";
		s_E353_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AC1";
		s_E354_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AC3";
		s_E355_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AC5";
		s_E356_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AC7";
		s_E357_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AC9";
		s_E358_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ACB";
		s_E359_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ACD";
		s_E360_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ACF";
		s_E361_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AD1";
		s_E362_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AD3";
		s_E363_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AD5";
		s_E364_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AD7";
		s_E365_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AD9";
		s_E366_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ADB";
		s_E367_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ADD";
		s_E368_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ADF";
		s_E369_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AE1";
		s_E370_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AE3";
		s_E371_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AE5";
		s_E372_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AE7";
		s_E373_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AE9";
		s_E374_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AEB";
		s_E375_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AED";
		s_E376_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AEF";
		s_E377_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AF1";
		s_E378_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AF3";
		s_E379_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AF5";
		s_E380_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AF7";
		s_E381_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AF9";
		s_E382_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AFB";
		s_E383_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AFD";
		s_E384_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"AFF";
		s_E385_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B01";
		s_E386_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B03";
		s_E387_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B05";
		s_E388_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B07";
		s_E389_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B09";
		s_E390_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B0B";
		s_E391_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B0D";
		s_E392_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B0F";
		s_E393_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B11";
		s_E394_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B13";
		s_E395_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B15";
		s_E396_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B17";
		s_E397_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B19";
		s_E398_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B1B";
		s_E399_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B1D";
		s_E400_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B1F";
		s_E401_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B21";
		s_E402_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B23";
		s_E403_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B25";
		s_E404_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B27";
		s_E405_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B29";
		s_E406_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B2B";
		s_E407_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B2D";
		s_E408_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B2F";
		s_E409_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B31";
		s_E410_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B33";
		s_E411_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B35";
		s_E412_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B37";
		s_E413_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B39";
		s_E414_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B3B";
		s_E415_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B3D";
		s_E416_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B3F";
		s_E417_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B41";
		s_E418_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B43";
		s_E419_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B45";
		s_E420_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B47";
		s_E421_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B49";
		s_E422_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B4B";
		s_E423_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B4D";
		s_E424_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B4F";
		s_E425_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B51";
		s_E426_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B53";
		s_E427_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B55";
		s_E428_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B57";
		s_E429_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B59";
		s_E430_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B5B";
		s_E431_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B5D";
		s_E432_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B5F";
		s_E433_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B61";
		s_E434_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B63";
		s_E435_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B65";
		s_E436_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B67";
		s_E437_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B69";
		s_E438_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B6B";
		s_E439_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B6D";
		s_E440_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B6F";
		s_E441_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B71";
		s_E442_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B73";
		s_E443_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B75";
		s_E444_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B77";
		s_E445_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B79";
		s_E446_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B7B";
		s_E447_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B7D";
		s_E448_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B7F";
		s_E449_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B81";
		s_E450_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B83";
		s_E451_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B85";
		s_E452_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B87";
		s_E453_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B89";
		s_E454_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B8B";
		s_E455_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B8D";
		s_E456_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B8F";
		s_E457_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B91";
		s_E458_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B93";
		s_E459_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B95";
		s_E460_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B97";
		s_E461_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B99";
		s_E462_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B9B";
		s_E463_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B9D";
		s_E464_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"B9F";
		s_E465_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BA1";
		s_E466_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BA3";
		s_E467_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BA5";
		s_E468_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BA7";
		s_E469_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BA9";
		s_E470_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BAB";
		s_E471_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BAD";
		s_E472_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BAF";
		s_E473_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BB1";
		s_E474_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BB3";
		s_E475_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BB5";
		s_E476_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BB7";
		s_E477_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BB9";
		s_E478_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BBB";
		s_E479_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BBD";
		s_E480_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BBF";
		s_E481_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BC1";
		s_E482_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BC3";
		s_E483_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BC5";
		s_E484_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BC7";
		s_E485_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BC9";
		s_E486_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BCB";
		s_E487_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BCD";
		s_E488_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BCF";
		s_E489_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BD1";
		s_E490_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BD3";
		s_E491_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BD5";
		s_E492_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BD7";
		s_E493_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BD9";
		s_E494_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BDB";
		s_E495_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BDD";
		s_E496_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BDF";
		s_E497_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BE1";
		s_E498_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BE3";
		s_E499_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BE5";
		s_E500_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BE7";
		s_E501_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BE9";
		s_E502_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BEB";
		s_E503_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BED";
		s_E504_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BEF";
		s_E505_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BF1";
		s_E506_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BF3";
		s_E507_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BF5";
		s_E508_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BF7";
		s_E509_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BF9";
		s_E510_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BFB";
		s_E511_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BFD";
		s_E512_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"BFF";
		s_E513_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C01";
		s_E514_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C03";
		s_E515_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C05";
		s_E516_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C07";
		s_E517_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C09";
		s_E518_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C0B";
		s_E519_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C0D";
		s_E520_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C0F";
		s_E521_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C11";
		s_E522_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C13";
		s_E523_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C15";
		s_E524_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C17";
		s_E525_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C19";
		s_E526_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C1B";
		s_E527_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C1D";
		s_E528_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C1F";
		s_E529_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C21";
		s_E530_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C23";
		s_E531_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C25";
		s_E532_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C27";
		s_E533_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C29";
		s_E534_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C2B";
		s_E535_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C2D";
		s_E536_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C2F";
		s_E537_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C31";
		s_E538_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C33";
		s_E539_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C35";
		s_E540_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C37";
		s_E541_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C39";
		s_E542_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C3B";
		s_E543_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C3D";
		s_E544_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C3F";
		s_E545_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C41";
		s_E546_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C43";
		s_E547_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C45";
		s_E548_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C47";
		s_E549_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C49";
		s_E550_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C4B";
		s_E551_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C4D";
		s_E552_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C4F";
		s_E553_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C51";
		s_E554_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C53";
		s_E555_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C55";
		s_E556_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C57";
		s_E557_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C59";
		s_E558_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C5B";
		s_E559_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C5D";
		s_E560_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C5F";
		s_E561_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C61";
		s_E562_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C63";
		s_E563_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C65";
		s_E564_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C67";
		s_E565_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C69";
		s_E566_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C6B";
		s_E567_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C6D";
		s_E568_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C6F";
		s_E569_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C71";
		s_E570_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C73";
		s_E571_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C75";
		s_E572_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C77";
		s_E573_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C79";
		s_E574_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C7B";
		s_E575_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C7D";
		s_E576_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C7F";
		s_E577_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C81";
		s_E578_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C83";
		s_E579_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C85";
		s_E580_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C87";
		s_E581_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C89";
		s_E582_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C8B";
		s_E583_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C8D";
		s_E584_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C8F";
		s_E585_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C91";
		s_E586_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C93";
		s_E587_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C95";
		s_E588_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C97";
		s_E589_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C99";
		s_E590_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C9B";
		s_E591_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C9D";
		s_E592_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"C9F";
		s_E593_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CA1";
		s_E594_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CA3";
		s_E595_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CA5";
		s_E596_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CA7";
		s_E597_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CA9";
		s_E598_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CAB";
		s_E599_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CAD";
		s_E600_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CAF";
		s_E601_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CB1";
		s_E602_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CB3";
		s_E603_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CB5";
		s_E604_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CB7";
		s_E605_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CB9";
		s_E606_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CBB";
		s_E607_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CBD";
		s_E608_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CBF";
		s_E609_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CC1";
		s_E610_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CC3";
		s_E611_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CC5";
		s_E612_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CC7";
		s_E613_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CC9";
		s_E614_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CCB";
		s_E615_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CCD";
		s_E616_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CCF";
		s_E617_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CD1";
		s_E618_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CD3";
		s_E619_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CD5";
		s_E620_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CD7";
		s_E621_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CD9";
		s_E622_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CDB";
		s_E623_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CDD";
		s_E624_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CDF";
		s_E625_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CE1";
		s_E626_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CE3";
		s_E627_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CE5";
		s_E628_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CE7";
		s_E629_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CE9";
		s_E630_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CEB";
		s_E631_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CED";
		s_E632_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CEF";
		s_E633_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CF1";
		s_E634_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CF3";
		s_E635_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CF5";
		s_E636_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CF7";
		s_E637_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CF9";
		s_E638_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CFB";
		s_E639_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CFD";
		s_E640_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"CFF";
		s_E641_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D01";
		s_E642_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D03";
		s_E643_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D05";
		s_E644_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D07";
		s_E645_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D09";
		s_E646_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D0B";
		s_E647_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D0D";
		s_E648_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D0F";
		s_E649_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D11";
		s_E650_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D13";
		s_E651_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D15";
		s_E652_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D17";
		s_E653_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D19";
		s_E654_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D1B";
		s_E655_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D1D";
		s_E656_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D1F";
		s_E657_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D21";
		s_E658_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D23";
		s_E659_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D25";
		s_E660_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D27";
		s_E661_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D29";
		s_E662_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D2B";
		s_E663_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D2D";
		s_E664_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D2F";
		s_E665_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D31";
		s_E666_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D33";
		s_E667_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D35";
		s_E668_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D37";
		s_E669_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D39";
		s_E670_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D3B";
		s_E671_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D3D";
		s_E672_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D3F";
		s_E673_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D41";
		s_E674_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D43";
		s_E675_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D45";
		s_E676_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D47";
		s_E677_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D49";
		s_E678_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D4B";
		s_E679_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D4D";
		s_E680_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D4F";
		s_E681_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D51";
		s_E682_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D53";
		s_E683_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D55";
		s_E684_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D57";
		s_E685_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D59";
		s_E686_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D5B";
		s_E687_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D5D";
		s_E688_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D5F";
		s_E689_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D61";
		s_E690_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D63";
		s_E691_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D65";
		s_E692_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D67";
		s_E693_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D69";
		s_E694_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D6B";
		s_E695_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D6D";
		s_E696_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D6F";
		s_E697_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D71";
		s_E698_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D73";
		s_E699_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D75";
		s_E700_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D77";
		s_E701_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D79";
		s_E702_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D7B";
		s_E703_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D7D";
		s_E704_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D7F";
		s_E705_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D81";
		s_E706_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D83";
		s_E707_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D85";
		s_E708_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D87";
		s_E709_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D89";
		s_E710_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D8B";
		s_E711_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D8D";
		s_E712_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D8F";
		s_E713_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D91";
		s_E714_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D93";
		s_E715_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D95";
		s_E716_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D97";
		s_E717_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D99";
		s_E718_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D9B";
		s_E719_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D9D";
		s_E720_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"D9F";
		s_E721_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DA1";
		s_E722_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DA3";
		s_E723_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DA5";
		s_E724_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DA7";
		s_E725_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DA9";
		s_E726_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DAB";
		s_E727_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DAD";
		s_E728_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DAF";
		s_E729_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DB1";
		s_E730_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DB3";
		s_E731_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DB5";
		s_E732_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DB7";
		s_E733_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DB9";
		s_E734_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DBB";
		s_E735_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DBD";
		s_E736_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DBF";
		s_E737_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DC1";
		s_E738_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DC3";
		s_E739_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DC5";
		s_E740_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DC7";
		s_E741_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DC9";
		s_E742_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DCB";
		s_E743_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DCD";
		s_E744_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DCF";
		s_E745_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DD1";
		s_E746_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DD3";
		s_E747_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DD5";
		s_E748_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DD7";
		s_E749_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DD9";
		s_E750_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DDB";
		s_E751_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DDD";
		s_E752_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DDF";
		s_E753_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DE1";
		s_E754_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DE3";
		s_E755_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DE5";
		s_E756_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DE7";
		s_E757_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DE9";
		s_E758_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DEB";
		s_E759_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DED";
		s_E760_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DEF";
		s_E761_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DF1";
		s_E762_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DF3";
		s_E763_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DF5";
		s_E764_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DF7";
		s_E765_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DF9";
		s_E766_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DFB";
		s_E767_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DFD";
		s_E768_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"DFF";
		s_E769_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E01";
		s_E770_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E03";
		s_E771_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E05";
		s_E772_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E07";
		s_E773_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E09";
		s_E774_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E0B";
		s_E775_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E0D";
		s_E776_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E0F";
		s_E777_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E11";
		s_E778_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E13";
		s_E779_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E15";
		s_E780_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E17";
		s_E781_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E19";
		s_E782_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E1B";
		s_E783_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E1D";
		s_E784_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E1F";
		s_E785_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E21";
		s_E786_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E23";
		s_E787_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E25";
		s_E788_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E27";
		s_E789_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E29";
		s_E790_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E2B";
		s_E791_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E2D";
		s_E792_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E2F";
		s_E793_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E31";
		s_E794_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E33";
		s_E795_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E35";
		s_E796_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E37";
		s_E797_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E39";
		s_E798_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E3B";
		s_E799_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E3D";
		s_E800_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E3F";
		s_E801_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E41";
		s_E802_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E43";
		s_E803_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E45";
		s_E804_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E47";
		s_E805_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E49";
		s_E806_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E4B";
		s_E807_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E4D";
		s_E808_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E4F";
		s_E809_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E51";
		s_E810_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E53";
		s_E811_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E55";
		s_E812_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E57";
		s_E813_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E59";
		s_E814_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E5B";
		s_E815_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E5D";
		s_E816_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E5F";
		s_E817_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E61";
		s_E818_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E63";
		s_E819_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E65";
		s_E820_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E67";
		s_E821_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E69";
		s_E822_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E6B";
		s_E823_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E6D";
		s_E824_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E6F";
		s_E825_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E71";
		s_E826_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E73";
		s_E827_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E75";
		s_E828_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E77";
		s_E829_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E79";
		s_E830_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E7B";
		s_E831_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E7D";
		s_E832_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E7F";
		s_E833_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E81";
		s_E834_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E83";
		s_E835_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E85";
		s_E836_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E87";
		s_E837_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E89";
		s_E838_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E8B";
		s_E839_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E8D";
		s_E840_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E8F";
		s_E841_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E91";
		s_E842_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E93";
		s_E843_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E95";
		s_E844_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E97";
		s_E845_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E99";
		s_E846_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E9B";
		s_E847_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E9D";
		s_E848_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"E9F";
		s_E849_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EA1";
		s_E850_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EA3";
		s_E851_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EA5";
		s_E852_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EA7";
		s_E853_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EA9";
		s_E854_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EAB";
		s_E855_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EAD";
		s_E856_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EAF";
		s_E857_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EB1";
		s_E858_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EB3";
		s_E859_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EB5";
		s_E860_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EB7";
		s_E861_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EB9";
		s_E862_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EBB";
		s_E863_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EBD";
		s_E864_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EBF";
		s_E865_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EC1";
		s_E866_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EC3";
		s_E867_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EC5";
		s_E868_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EC7";
		s_E869_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EC9";
		s_E870_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ECB";
		s_E871_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ECD";
		s_E872_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ECF";
		s_E873_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ED1";
		s_E874_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ED3";
		s_E875_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ED5";
		s_E876_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ED7";
		s_E877_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"ED9";
		s_E878_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EDB";
		s_E879_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EDD";
		s_E880_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EDF";
		s_E881_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EE1";
		s_E882_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EE3";
		s_E883_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EE5";
		s_E884_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EE7";
		s_E885_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EE9";
		s_E886_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EEB";
		s_E887_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EED";
		s_E888_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EEF";
		s_E889_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EF1";
		s_E890_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EF3";
		s_E891_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EF5";
		s_E892_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EF7";
		s_E893_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EF9";
		s_E894_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EFB";
		s_E895_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EFD";
		s_E896_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"EFF";
		s_E897_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F01";
		s_E898_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F03";
		s_E899_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F05";
		s_E900_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F07";
		s_E901_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F09";
		s_E902_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F0B";
		s_E903_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F0D";
		s_E904_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F0F";
		s_E905_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F11";
		s_E906_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F13";
		s_E907_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F15";
		s_E908_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F17";
		s_E909_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F19";
		s_E910_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F1B";
		s_E911_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F1D";
		s_E912_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F1F";
		s_E913_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F21";
		s_E914_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F23";
		s_E915_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F25";
		s_E916_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F27";
		s_E917_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F29";
		s_E918_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F2B";
		s_E919_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F2D";
		s_E920_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F2F";
		s_E921_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F31";
		s_E922_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F33";
		s_E923_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F35";
		s_E924_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F37";
		s_E925_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F39";
		s_E926_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F3B";
		s_E927_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F3D";
		s_E928_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F3F";
		s_E929_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F41";
		s_E930_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F43";
		s_E931_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F45";
		s_E932_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F47";
		s_E933_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F49";
		s_E934_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F4B";
		s_E935_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F4D";
		s_E936_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F4F";
		s_E937_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F51";
		s_E938_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F53";
		s_E939_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F55";
		s_E940_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F57";
		s_E941_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F59";
		s_E942_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F5B";
		s_E943_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F5D";
		s_E944_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F5F";
		s_E945_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F61";
		s_E946_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F63";
		s_E947_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F65";
		s_E948_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F67";
		s_E949_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F69";
		s_E950_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F6B";
		s_E951_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F6D";
		s_E952_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F6F";
		s_E953_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F71";
		s_E954_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F73";
		s_E955_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F75";
		s_E956_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F77";
		s_E957_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F79";
		s_E958_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F7B";
		s_E959_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F7D";
		s_E960_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F7F";
		s_E961_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F81";
		s_E962_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F83";
		s_E963_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F85";
		s_E964_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F87";
		s_E965_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F89";
		s_E966_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F8B";
		s_E967_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F8D";
		s_E968_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F8F";
		s_E969_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F91";
		s_E970_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F93";
		s_E971_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F95";
		s_E972_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F97";
		s_E973_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F99";
		s_E974_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F9B";
		s_E975_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F9D";
		s_E976_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"F9F";
		s_E977_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FA1";
		s_E978_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FA3";
		s_E979_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FA5";
		s_E980_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FA7";
		s_E981_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FA9";
		s_E982_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FAB";
		s_E983_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FAD";
		s_E984_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FAF";
		s_E985_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FB1";
		s_E986_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FB3";
		s_E987_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FB5";
		s_E988_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FB7";
		s_E989_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FB9";
		s_E990_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FBB";
		s_E991_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FBD";
		s_E992_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FBF";
		s_E993_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FC1";
		s_E994_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FC3";
		s_E995_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FC5";
		s_E996_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FC7";
		s_E997_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FC9";
		s_E998_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FCB";
		s_E999_C1_H_Pos			  :std_logic_vector(11 downto 0) := x"FCD";
		s_E1000_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FCF";
		s_E1001_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FD1";
		s_E1002_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FD3";
		s_E1003_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FD5";
		s_E1004_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FD7";
		s_E1005_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FD9";
		s_E1006_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FDB";
		s_E1007_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FDD";
		s_E1008_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FDF";
		s_E1009_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FE1";
		s_E1010_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FE3";
		s_E1011_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FE5";
		s_E1012_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FE7";
		s_E1013_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FE9";
		s_E1014_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FEB";
		s_E1015_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FED";
		s_E1016_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FEF";
		s_E1017_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FF1";
		s_E1018_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FF3";
		s_E1019_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FF5";
		s_E1020_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FF7";
		s_E1021_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FF9";
		s_E1022_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FFB";
		s_E1023_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FFD";
		s_E1024_C1_H_Pos		  :std_logic_vector(11 downto 0) := x"FFF";

		s_E2_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"801";
		s_E3_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"803";
		s_E4_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"805";
		s_E5_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"807";
		s_E6_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"809";
		s_E7_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"80B";
		s_E8_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"80D";
		s_E9_C1_L_Pos        	  :std_logic_vector(11 downto 0) := x"80F";
		s_E10_C1_L_Pos       	  :std_logic_vector(11 downto 0) := x"811";
		s_E11_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"813";
		s_E12_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"815";
		s_E13_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"817";
		s_E14_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"819";
		s_E15_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"81B";
		s_E16_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"81D";
		s_E17_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"81F";
		s_E18_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"821";
		s_E19_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"823";
		s_E20_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"825";
		s_E21_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"827";
		s_E22_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"829";
		s_E23_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"82B";
		s_E24_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"82D";
		s_E25_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"82F";
		s_E26_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"831";
		s_E27_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"833";
		s_E28_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"835";
		s_E29_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"837";
		s_E30_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"839";
		s_E31_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"83B";
		s_E32_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"83D";
		s_E33_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"83F";
		s_E34_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"841";
		s_E35_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"843";
		s_E36_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"845";
		s_E37_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"847";
		s_E38_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"849";
		s_E39_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"84B";
		s_E40_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"84D";
		s_E41_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"84F";
		s_E42_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"851";
		s_E43_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"853";
		s_E44_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"855";
		s_E45_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"857";
		s_E46_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"859";
		s_E47_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"85B";
		s_E48_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"85D";
		s_E49_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"85F";
		s_E50_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"861";
		s_E51_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"863";
		s_E52_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"865";
		s_E53_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"867";
		s_E54_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"869";
		s_E55_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"86B";
		s_E56_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"86D";
		s_E57_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"86F";
		s_E58_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"871";
		s_E59_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"873";
		s_E60_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"875";
		s_E61_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"877";
		s_E62_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"879";
		s_E63_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"87B";
		s_E64_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"87D";
		s_E65_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"87F";
		s_E66_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"881";
		s_E67_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"883";
		s_E68_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"885";
		s_E69_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"887";
		s_E70_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"889";
		s_E71_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"88B";
		s_E72_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"88D";
		s_E73_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"88F";
		s_E74_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"891";
		s_E75_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"893";
		s_E76_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"895";
		s_E77_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"897";
		s_E78_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"899";
		s_E79_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"89B";
		s_E80_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"89D";
		s_E81_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"89F";
		s_E82_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8A1";
		s_E83_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8A3";
		s_E84_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8A5";
		s_E85_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8A7";
		s_E86_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8A9";
		s_E87_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8AB";
		s_E88_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8AD";
		s_E89_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8AF";
		s_E90_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8B1";
		s_E91_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8B3";
		s_E92_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8B5";
		s_E93_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8B7";
		s_E94_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8B9";
		s_E95_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8BB";
		s_E96_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8BD";
		s_E97_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8BF";
		s_E98_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8C1";
		s_E99_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8C3";
		s_E100_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8C5";
		s_E101_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8C7";
		s_E102_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8C9";
		s_E103_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8CB";
		s_E104_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8CD";
		s_E105_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8CF";
		s_E106_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8D1";
		s_E107_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8D3";
		s_E108_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8D5";
		s_E109_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8D7";
		s_E110_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8D9";
		s_E111_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8DB";
		s_E112_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8DD";
		s_E113_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8DF";
		s_E114_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8E1";
		s_E115_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8E3";
		s_E116_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8E5";
		s_E117_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8E7";
		s_E118_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8E9";
		s_E119_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8EB";
		s_E120_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8ED";
		s_E121_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8EF";
		s_E122_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8F1";
		s_E123_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8F3";
		s_E124_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8F5";
		s_E125_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8F7";
		s_E126_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8F9";
		s_E127_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8FB";
		s_E128_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8FD";
		s_E129_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"8FF";
		s_E130_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"901";
		s_E131_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"903";
		s_E132_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"905";
		s_E133_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"907";
		s_E134_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"909";
		s_E135_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"90B";
		s_E136_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"90D";
		s_E137_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"90F";
		s_E138_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"911";
		s_E139_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"913";
		s_E140_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"915";
		s_E141_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"917";
		s_E142_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"919";
		s_E143_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"91B";
		s_E144_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"91D";
		s_E145_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"91F";
		s_E146_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"921";
		s_E147_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"923";
		s_E148_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"925";
		s_E149_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"927";
		s_E150_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"929";
		s_E151_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"92B";
		s_E152_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"92D";
		s_E153_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"92F";
		s_E154_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"931";
		s_E155_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"933";
		s_E156_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"935";
		s_E157_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"937";
		s_E158_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"939";
		s_E159_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"93B";
		s_E160_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"93D";
		s_E161_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"93F";
		s_E162_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"941";
		s_E163_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"943";
		s_E164_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"945";
		s_E165_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"947";
		s_E166_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"949";
		s_E167_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"94B";
		s_E168_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"94D";
		s_E169_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"94F";
		s_E170_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"951";
		s_E171_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"953";
		s_E172_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"955";
		s_E173_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"957";
		s_E174_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"959";
		s_E175_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"95B";
		s_E176_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"95D";
		s_E177_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"95F";
		s_E178_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"961";
		s_E179_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"963";
		s_E180_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"965";
		s_E181_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"967";
		s_E182_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"969";
		s_E183_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"96B";
		s_E184_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"96D";
		s_E185_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"96F";
		s_E186_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"971";
		s_E187_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"973";
		s_E188_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"975";
		s_E189_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"977";
		s_E190_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"979";
		s_E191_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"97B";
		s_E192_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"97D";
		s_E193_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"97F";
		s_E194_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"981";
		s_E195_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"983";
		s_E196_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"985";
		s_E197_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"987";
		s_E198_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"989";
		s_E199_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"98B";
		s_E200_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"98D";
		s_E201_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"98F";
		s_E202_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"991";
		s_E203_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"993";
		s_E204_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"995";
		s_E205_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"997";
		s_E206_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"999";
		s_E207_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"99B";
		s_E208_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"99D";
		s_E209_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"99F";
		s_E210_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9A1";
		s_E211_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9A3";
		s_E212_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9A5";
		s_E213_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9A7";
		s_E214_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9A9";
		s_E215_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9AB";
		s_E216_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9AD";
		s_E217_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9AF";
		s_E218_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9B1";
		s_E219_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9B3";
		s_E220_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9B5";
		s_E221_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9B7";
		s_E222_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9B9";
		s_E223_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9BB";
		s_E224_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9BD";
		s_E225_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9BF";
		s_E226_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9C1";
		s_E227_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9C3";
		s_E228_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9C5";
		s_E229_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9C7";
		s_E230_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9C9";
		s_E231_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9CB";
		s_E232_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9CD";
		s_E233_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9CF";
		s_E234_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9D1";
		s_E235_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9D3";
		s_E236_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9D5";
		s_E237_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9D7";
		s_E238_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9D9";
		s_E239_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9DB";
		s_E240_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9DD";
		s_E241_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9DF";
		s_E242_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9E1";
		s_E243_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9E3";
		s_E244_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9E5";
		s_E245_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9E7";
		s_E246_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9E9";
		s_E247_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9EB";
		s_E248_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9ED";
		s_E249_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9EF";
		s_E250_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9F1";
		s_E251_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9F3";
		s_E252_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9F5";
		s_E253_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9F7";
		s_E254_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9F9";
		s_E255_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9FB";
		s_E256_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9FD";
		s_E257_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"9FF";
		s_E258_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A01";
		s_E259_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A03";
		s_E260_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A05";
		s_E261_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A07";
		s_E262_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A09";
		s_E263_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A0B";
		s_E264_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A0D";
		s_E265_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A0F";
		s_E266_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A11";
		s_E267_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A13";
		s_E268_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A15";
		s_E269_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A17";
		s_E270_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A19";
		s_E271_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A1B";
		s_E272_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A1D";
		s_E273_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A1F";
		s_E274_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A21";
		s_E275_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A23";
		s_E276_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A25";
		s_E277_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A27";
		s_E278_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A29";
		s_E279_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A2B";
		s_E280_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A2D";
		s_E281_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A2F";
		s_E282_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A31";
		s_E283_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A33";
		s_E284_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A35";
		s_E285_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A37";
		s_E286_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A39";
		s_E287_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A3B";
		s_E288_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A3D";
		s_E289_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A3F";
		s_E290_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A41";
		s_E291_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A43";
		s_E292_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A45";
		s_E293_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A47";
		s_E294_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A49";
		s_E295_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A4B";
		s_E296_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A4D";
		s_E297_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A4F";
		s_E298_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A51";
		s_E299_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A53";
		s_E300_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A55";
		s_E301_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A57";
		s_E302_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A59";
		s_E303_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A5B";
		s_E304_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A5D";
		s_E305_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A5F";
		s_E306_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A61";
		s_E307_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A63";
		s_E308_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A65";
		s_E309_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A67";
		s_E310_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A69";
		s_E311_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A6B";
		s_E312_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A6D";
		s_E313_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A6F";
		s_E314_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A71";
		s_E315_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A73";
		s_E316_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A75";
		s_E317_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A77";
		s_E318_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A79";
		s_E319_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A7B";
		s_E320_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A7D";
		s_E321_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A7F";
		s_E322_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A81";
		s_E323_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A83";
		s_E324_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A85";
		s_E325_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A87";
		s_E326_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A89";
		s_E327_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A8B";
		s_E328_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A8D";
		s_E329_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A8F";
		s_E330_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A91";
		s_E331_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A93";
		s_E332_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A95";
		s_E333_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A97";
		s_E334_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A99";
		s_E335_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A9B";
		s_E336_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A9D";
		s_E337_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"A9F";
		s_E338_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AA1";
		s_E339_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AA3";
		s_E340_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AA5";
		s_E341_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AA7";
		s_E342_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AA9";
		s_E343_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AAB";
		s_E344_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AAD";
		s_E345_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AAF";
		s_E346_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AB1";
		s_E347_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AB3";
		s_E348_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AB5";
		s_E349_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AB7";
		s_E350_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AB9";
		s_E351_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ABB";
		s_E352_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ABD";
		s_E353_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ABF";
		s_E354_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AC1";
		s_E355_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AC3";
		s_E356_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AC5";
		s_E357_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AC7";
		s_E358_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AC9";
		s_E359_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ACB";
		s_E360_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ACD";
		s_E361_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ACF";
		s_E362_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AD1";
		s_E363_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AD3";
		s_E364_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AD5";
		s_E365_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AD7";
		s_E366_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AD9";
		s_E367_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ADB";
		s_E368_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ADD";
		s_E369_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ADF";
		s_E370_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AE1";
		s_E371_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AE3";
		s_E372_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AE5";
		s_E373_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AE7";
		s_E374_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AE9";
		s_E375_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AEB";
		s_E376_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AED";
		s_E377_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AEF";
		s_E378_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AF1";
		s_E379_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AF3";
		s_E380_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AF5";
		s_E381_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AF7";
		s_E382_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AF9";
		s_E383_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AFB";
		s_E384_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AFD";
		s_E385_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"AFF";
		s_E386_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B01";
		s_E387_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B03";
		s_E388_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B05";
		s_E389_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B07";
		s_E390_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B09";
		s_E391_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B0B";
		s_E392_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B0D";
		s_E393_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B0F";
		s_E394_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B11";
		s_E395_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B13";
		s_E396_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B15";
		s_E397_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B17";
		s_E398_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B19";
		s_E399_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B1B";
		s_E400_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B1D";
		s_E401_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B1F";
		s_E402_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B21";
		s_E403_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B23";
		s_E404_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B25";
		s_E405_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B27";
		s_E406_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B29";
		s_E407_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B2B";
		s_E408_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B2D";
		s_E409_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B2F";
		s_E410_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B31";
		s_E411_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B33";
		s_E412_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B35";
		s_E413_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B37";
		s_E414_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B39";
		s_E415_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B3B";
		s_E416_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B3D";
		s_E417_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B3F";
		s_E418_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B41";
		s_E419_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B43";
		s_E420_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B45";
		s_E421_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B47";
		s_E422_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B49";
		s_E423_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B4B";
		s_E424_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B4D";
		s_E425_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B4F";
		s_E426_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B51";
		s_E427_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B53";
		s_E428_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B55";
		s_E429_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B57";
		s_E430_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B59";
		s_E431_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B5B";
		s_E432_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B5D";
		s_E433_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B5F";
		s_E434_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B61";
		s_E435_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B63";
		s_E436_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B65";
		s_E437_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B67";
		s_E438_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B69";
		s_E439_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B6B";
		s_E440_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B6D";
		s_E441_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B6F";
		s_E442_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B71";
		s_E443_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B73";
		s_E444_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B75";
		s_E445_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B77";
		s_E446_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B79";
		s_E447_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B7B";
		s_E448_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B7D";
		s_E449_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B7F";
		s_E450_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B81";
		s_E451_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B83";
		s_E452_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B85";
		s_E453_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B87";
		s_E454_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B89";
		s_E455_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B8B";
		s_E456_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B8D";
		s_E457_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B8F";
		s_E458_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B91";
		s_E459_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B93";
		s_E460_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B95";
		s_E461_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B97";
		s_E462_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B99";
		s_E463_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B9B";
		s_E464_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B9D";
		s_E465_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"B9F";
		s_E466_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BA1";
		s_E467_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BA3";
		s_E468_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BA5";
		s_E469_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BA7";
		s_E470_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BA9";
		s_E471_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BAB";
		s_E472_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BAD";
		s_E473_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BAF";
		s_E474_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BB1";
		s_E475_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BB3";
		s_E476_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BB5";
		s_E477_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BB7";
		s_E478_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BB9";
		s_E479_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BBB";
		s_E480_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BBD";
		s_E481_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BBF";
		s_E482_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BC1";
		s_E483_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BC3";
		s_E484_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BC5";
		s_E485_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BC7";
		s_E486_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BC9";
		s_E487_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BCB";
		s_E488_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BCD";
		s_E489_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BCF";
		s_E490_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BD1";
		s_E491_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BD3";
		s_E492_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BD5";
		s_E493_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BD7";
		s_E494_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BD9";
		s_E495_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BDB";
		s_E496_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BDD";
		s_E497_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BDF";
		s_E498_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BE1";
		s_E499_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BE3";
		s_E500_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BE5";
		s_E501_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BE7";
		s_E502_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BE9";
		s_E503_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BEB";
		s_E504_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BED";
		s_E505_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BEF";
		s_E506_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BF1";
		s_E507_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BF3";
		s_E508_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BF5";
		s_E509_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BF7";
		s_E510_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BF9";
		s_E511_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BFB";
		s_E512_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BFD";
		s_E513_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"BFF";
		s_E514_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C01";
		s_E515_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C03";
		s_E516_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C05";
		s_E517_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C07";
		s_E518_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C09";
		s_E519_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C0B";
		s_E520_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C0D";
		s_E521_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C0F";
		s_E522_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C11";
		s_E523_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C13";
		s_E524_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C15";
		s_E525_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C17";
		s_E526_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C19";
		s_E527_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C1B";
		s_E528_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C1D";
		s_E529_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C1F";
		s_E530_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C21";
		s_E531_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C23";
		s_E532_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C25";
		s_E533_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C27";
		s_E534_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C29";
		s_E535_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C2B";
		s_E536_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C2D";
		s_E537_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C2F";
		s_E538_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C31";
		s_E539_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C33";
		s_E540_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C35";
		s_E541_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C37";
		s_E542_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C39";
		s_E543_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C3B";
		s_E544_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C3D";
		s_E545_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C3F";
		s_E546_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C41";
		s_E547_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C43";
		s_E548_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C45";
		s_E549_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C47";
		s_E550_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C49";
		s_E551_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C4B";
		s_E552_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C4D";
		s_E553_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C4F";
		s_E554_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C51";
		s_E555_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C53";
		s_E556_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C55";
		s_E557_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C57";
		s_E558_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C59";
		s_E559_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C5B";
		s_E560_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C5D";
		s_E561_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C5F";
		s_E562_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C61";
		s_E563_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C63";
		s_E564_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C65";
		s_E565_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C67";
		s_E566_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C69";
		s_E567_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C6B";
		s_E568_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C6D";
		s_E569_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C6F";
		s_E570_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C71";
		s_E571_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C73";
		s_E572_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C75";
		s_E573_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C77";
		s_E574_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C79";
		s_E575_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C7B";
		s_E576_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C7D";
		s_E577_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C7F";
		s_E578_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C81";
		s_E579_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C83";
		s_E580_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C85";
		s_E581_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C87";
		s_E582_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C89";
		s_E583_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C8B";
		s_E584_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C8D";
		s_E585_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C8F";
		s_E586_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C91";
		s_E587_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C93";
		s_E588_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C95";
		s_E589_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C97";
		s_E590_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C99";
		s_E591_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C9B";
		s_E592_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C9D";
		s_E593_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"C9F";
		s_E594_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CA1";
		s_E595_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CA3";
		s_E596_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CA5";
		s_E597_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CA7";
		s_E598_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CA9";
		s_E599_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CAB";
		s_E600_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CAD";
		s_E601_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CAF";
		s_E602_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CB1";
		s_E603_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CB3";
		s_E604_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CB5";
		s_E605_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CB7";
		s_E606_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CB9";
		s_E607_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CBB";
		s_E608_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CBD";
		s_E609_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CBF";
		s_E610_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CC1";
		s_E611_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CC3";
		s_E612_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CC5";
		s_E613_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CC7";
		s_E614_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CC9";
		s_E615_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CCB";
		s_E616_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CCD";
		s_E617_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CCF";
		s_E618_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CD1";
		s_E619_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CD3";
		s_E620_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CD5";
		s_E621_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CD7";
		s_E622_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CD9";
		s_E623_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CDB";
		s_E624_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CDD";
		s_E625_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CDF";
		s_E626_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CE1";
		s_E627_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CE3";
		s_E628_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CE5";
		s_E629_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CE7";
		s_E630_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CE9";
		s_E631_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CEB";
		s_E632_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CED";
		s_E633_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CEF";
		s_E634_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CF1";
		s_E635_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CF3";
		s_E636_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CF5";
		s_E637_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CF7";
		s_E638_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CF9";
		s_E639_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CFB";
		s_E640_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CFD";
		s_E641_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"CFF";
		s_E642_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D01";
		s_E643_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D03";
		s_E644_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D05";
		s_E645_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D07";
		s_E646_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D09";
		s_E647_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D0B";
		s_E648_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D0D";
		s_E649_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D0F";
		s_E650_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D11";
		s_E651_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D13";
		s_E652_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D15";
		s_E653_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D17";
		s_E654_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D19";
		s_E655_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D1B";
		s_E656_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D1D";
		s_E657_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D1F";
		s_E658_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D21";
		s_E659_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D23";
		s_E660_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D25";
		s_E661_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D27";
		s_E662_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D29";
		s_E663_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D2B";
		s_E664_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D2D";
		s_E665_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D2F";
		s_E666_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D31";
		s_E667_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D33";
		s_E668_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D35";
		s_E669_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D37";
		s_E670_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D39";
		s_E671_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D3B";
		s_E672_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D3D";
		s_E673_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D3F";
		s_E674_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D41";
		s_E675_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D43";
		s_E676_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D45";
		s_E677_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D47";
		s_E678_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D49";
		s_E679_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D4B";
		s_E680_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D4D";
		s_E681_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D4F";
		s_E682_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D51";
		s_E683_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D53";
		s_E684_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D55";
		s_E685_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D57";
		s_E686_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D59";
		s_E687_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D5B";
		s_E688_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D5D";
		s_E689_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D5F";
		s_E690_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D61";
		s_E691_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D63";
		s_E692_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D65";
		s_E693_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D67";
		s_E694_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D69";
		s_E695_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D6B";
		s_E696_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D6D";
		s_E697_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D6F";
		s_E698_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D71";
		s_E699_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D73";
		s_E700_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D75";
		s_E701_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D77";
		s_E702_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D79";
		s_E703_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D7B";
		s_E704_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D7D";
		s_E705_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D7F";
		s_E706_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D81";
		s_E707_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D83";
		s_E708_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D85";
		s_E709_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D87";
		s_E710_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D89";
		s_E711_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D8B";
		s_E712_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D8D";
		s_E713_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D8F";
		s_E714_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D91";
		s_E715_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D93";
		s_E716_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D95";
		s_E717_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D97";
		s_E718_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D99";
		s_E719_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D9B";
		s_E720_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D9D";
		s_E721_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"D9F";
		s_E722_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DA1";
		s_E723_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DA3";
		s_E724_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DA5";
		s_E725_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DA7";
		s_E726_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DA9";
		s_E727_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DAB";
		s_E728_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DAD";
		s_E729_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DAF";
		s_E730_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DB1";
		s_E731_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DB3";
		s_E732_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DB5";
		s_E733_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DB7";
		s_E734_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DB9";
		s_E735_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DBB";
		s_E736_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DBD";
		s_E737_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DBF";
		s_E738_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DC1";
		s_E739_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DC3";
		s_E740_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DC5";
		s_E741_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DC7";
		s_E742_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DC9";
		s_E743_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DCB";
		s_E744_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DCD";
		s_E745_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DCF";
		s_E746_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DD1";
		s_E747_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DD3";
		s_E748_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DD5";
		s_E749_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DD7";
		s_E750_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DD9";
		s_E751_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DDB";
		s_E752_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DDD";
		s_E753_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DDF";
		s_E754_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DE1";
		s_E755_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DE3";
		s_E756_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DE5";
		s_E757_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DE7";
		s_E758_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DE9";
		s_E759_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DEB";
		s_E760_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DED";
		s_E761_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DEF";
		s_E762_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DF1";
		s_E763_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DF3";
		s_E764_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DF5";
		s_E765_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DF7";
		s_E766_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DF9";
		s_E767_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DFB";
		s_E768_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DFD";
		s_E769_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"DFF";
		s_E770_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E01";
		s_E771_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E03";
		s_E772_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E05";
		s_E773_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E07";
		s_E774_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E09";
		s_E775_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E0B";
		s_E776_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E0D";
		s_E777_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E0F";
		s_E778_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E11";
		s_E779_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E13";
		s_E780_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E15";
		s_E781_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E17";
		s_E782_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E19";
		s_E783_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E1B";
		s_E784_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E1D";
		s_E785_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E1F";
		s_E786_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E21";
		s_E787_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E23";
		s_E788_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E25";
		s_E789_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E27";
		s_E790_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E29";
		s_E791_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E2B";
		s_E792_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E2D";
		s_E793_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E2F";
		s_E794_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E31";
		s_E795_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E33";
		s_E796_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E35";
		s_E797_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E37";
		s_E798_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E39";
		s_E799_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E3B";
		s_E800_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E3D";
		s_E801_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E3F";
		s_E802_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E41";
		s_E803_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E43";
		s_E804_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E45";
		s_E805_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E47";
		s_E806_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E49";
		s_E807_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E4B";
		s_E808_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E4D";
		s_E809_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E4F";
		s_E810_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E51";
		s_E811_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E53";
		s_E812_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E55";
		s_E813_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E57";
		s_E814_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E59";
		s_E815_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E5B";
		s_E816_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E5D";
		s_E817_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E5F";
		s_E818_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E61";
		s_E819_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E63";
		s_E820_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E65";
		s_E821_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E67";
		s_E822_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E69";
		s_E823_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E6B";
		s_E824_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E6D";
		s_E825_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E6F";
		s_E826_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E71";
		s_E827_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E73";
		s_E828_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E75";
		s_E829_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E77";
		s_E830_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E79";
		s_E831_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E7B";
		s_E832_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E7D";
		s_E833_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E7F";
		s_E834_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E81";
		s_E835_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E83";
		s_E836_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E85";
		s_E837_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E87";
		s_E838_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E89";
		s_E839_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E8B";
		s_E840_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E8D";
		s_E841_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E8F";
		s_E842_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E91";
		s_E843_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E93";
		s_E844_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E95";
		s_E845_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E97";
		s_E846_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E99";
		s_E847_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E9B";
		s_E848_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E9D";
		s_E849_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"E9F";
		s_E850_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EA1";
		s_E851_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EA3";
		s_E852_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EA5";
		s_E853_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EA7";
		s_E854_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EA9";
		s_E855_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EAB";
		s_E856_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EAD";
		s_E857_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EAF";
		s_E858_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EB1";
		s_E859_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EB3";
		s_E860_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EB5";
		s_E861_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EB7";
		s_E862_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EB9";
		s_E863_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EBB";
		s_E864_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EBD";
		s_E865_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EBF";
		s_E866_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EC1";
		s_E867_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EC3";
		s_E868_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EC5";
		s_E869_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EC7";
		s_E870_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EC9";
		s_E871_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ECB";
		s_E872_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ECD";
		s_E873_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ECF";
		s_E874_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ED1";
		s_E875_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ED3";
		s_E876_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ED5";
		s_E877_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ED7";
		s_E878_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"ED9";
		s_E879_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EDB";
		s_E880_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EDD";
		s_E881_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EDF";
		s_E882_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EE1";
		s_E883_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EE3";
		s_E884_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EE5";
		s_E885_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EE7";
		s_E886_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EE9";
		s_E887_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EEB";
		s_E888_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EED";
		s_E889_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EEF";
		s_E890_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EF1";
		s_E891_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EF3";
		s_E892_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EF5";
		s_E893_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EF7";
		s_E894_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EF9";
		s_E895_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EFB";
		s_E896_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EFD";
		s_E897_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"EFF";
		s_E898_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F01";
		s_E899_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F03";
		s_E900_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F05";
		s_E901_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F07";
		s_E902_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F09";
		s_E903_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F0B";
		s_E904_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F0D";
		s_E905_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F0F";
		s_E906_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F11";
		s_E907_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F13";
		s_E908_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F15";
		s_E909_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F17";
		s_E910_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F19";
		s_E911_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F1B";
		s_E912_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F1D";
		s_E913_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F1F";
		s_E914_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F21";
		s_E915_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F23";
		s_E916_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F25";
		s_E917_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F27";
		s_E918_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F29";
		s_E919_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F2B";
		s_E920_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F2D";
		s_E921_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F2F";
		s_E922_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F31";
		s_E923_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F33";
		s_E924_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F35";
		s_E925_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F37";
		s_E926_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F39";
		s_E927_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F3B";
		s_E928_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F3D";
		s_E929_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F3F";
		s_E930_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F41";
		s_E931_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F43";
		s_E932_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F45";
		s_E933_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F47";
		s_E934_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F49";
		s_E935_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F4B";
		s_E936_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F4D";
		s_E937_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F4F";
		s_E938_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F51";
		s_E939_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F53";
		s_E940_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F55";
		s_E941_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F57";
		s_E942_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F59";
		s_E943_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F5B";
		s_E944_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F5D";
		s_E945_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F5F";
		s_E946_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F61";
		s_E947_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F63";
		s_E948_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F65";
		s_E949_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F67";
		s_E950_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F69";
		s_E951_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F6B";
		s_E952_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F6D";
		s_E953_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F6F";
		s_E954_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F71";
		s_E955_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F73";
		s_E956_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F75";
		s_E957_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F77";
		s_E958_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F79";
		s_E959_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F7B";
		s_E960_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F7D";
		s_E961_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F7F";
		s_E962_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F81";
		s_E963_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F83";
		s_E964_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F85";
		s_E965_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F87";
		s_E966_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F89";
		s_E967_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F8B";
		s_E968_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F8D";
		s_E969_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F8F";
		s_E970_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F91";
		s_E971_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F93";
		s_E972_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F95";
		s_E973_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F97";
		s_E974_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F99";
		s_E975_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F9B";
		s_E976_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F9D";
		s_E977_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"F9F";
		s_E978_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FA1";
		s_E979_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FA3";
		s_E980_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FA5";
		s_E981_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FA7";
		s_E982_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FA9";
		s_E983_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FAB";
		s_E984_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FAD";
		s_E985_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FAF";
		s_E986_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FB1";
		s_E987_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FB3";
		s_E988_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FB5";
		s_E989_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FB7";
		s_E990_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FB9";
		s_E991_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FBB";
		s_E992_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FBD";
		s_E993_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FBF";
		s_E994_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FC1";
		s_E995_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FC3";
		s_E996_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FC5";
		s_E997_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FC7";
		s_E998_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FC9";
		s_E999_C1_L_Pos			  :std_logic_vector(11 downto 0) := x"FCB";
		s_E1000_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FCD";
		s_E1001_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FCF";
		s_E1002_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FD1";
		s_E1003_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FD3";
		s_E1004_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FD5";
		s_E1005_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FD7";
		s_E1006_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FD9";
		s_E1007_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FDB";
		s_E1008_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FDD";
		s_E1009_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FDF";
		s_E1010_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FE1";
		s_E1011_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FE3";
		s_E1012_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FE5";
		s_E1013_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FE7";
		s_E1014_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FE9";
		s_E1015_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FEB";
		s_E1016_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FED";
		s_E1017_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FEF";
		s_E1018_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FF1";
		s_E1019_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FF3";
		s_E1020_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FF5";
		s_E1021_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FF7";
		s_E1022_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FF9";
		s_E1023_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FFB";
		s_E1024_C1_L_Pos		  :std_logic_vector(11 downto 0) := x"FFD"


		

      );

  --+----------
  -- Port name declarations
  --+----------
 port   (
       CLK100     			   :in  std_logic;
       RST        			   :in  std_logic;
       
       DATA1                   :in  std_logic_vector(WdVecSize_g-5 downto 0);
       DATARDY1                :in  std_logic;
       DATA2                   :in  std_logic_vector(WdVecSize_g-5 downto 0);
       DATARDY2                :in  std_logic;
        
--       THRESHOLD  :in  std_logic_vector(NibbleSize_g-1 downto 0);
       
	   ADD_TIMP_FLAG 		   :out std_logic;
	   ADD_TIMP_FLAG_pos 	   :out std_logic;
	   
	   o_DATA_OUT_C1  		   :out std_logic_vector(11 downto 0);
	   o_DATA_OUT_C2  		   :out std_logic_vector(11 downto 0);
							   
       i_PEAK_THD          	   :in std_logic_vector(11 downto 0);
       i_PEAK_THD_pos          :in std_logic_vector(11 downto 0);

	   o_Energy_Bin_1    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_2    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_3    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_4    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_5    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_6    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_7    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_8    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_9    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_10   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_11   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_12   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_13   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_14   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_15   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_16   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_17   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_18   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_19   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_20   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_21   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_22   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_23   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_24   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_25   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_26   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_27   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_28   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_29   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_30   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_31   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_32   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_33   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_34   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_35   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_36   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_37   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_38   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_39   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_40   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_41   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_42   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_43   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_44   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_45   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_46   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_47   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_48   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_49   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_50   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_51   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_52   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_53   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_54   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_55   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_56   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_57   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_58   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_59   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_60   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_61   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_62   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_63   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_64   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_65   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_66   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_67   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_68   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_69   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_70   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_71   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_72   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_73   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_74   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_75   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_76   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_77   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_78   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_79   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_80   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_81   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_82   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_83   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_84   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_85   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_86   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_87   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_88   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_89   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_90   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_91   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_92   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_93   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_94   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_95   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_96   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_97   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_98   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_99   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_100  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_101  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_102  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_103  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_104  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_105  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_106  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_107  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_108  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_109  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_110  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_111  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_112  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_113  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_114  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_115  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_116  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_117  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_118  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_119  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_120  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_121  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_122  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_123  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_124  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_125  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_126  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_127  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_128  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_129  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_130  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_131  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_132  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_133  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_134  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_135  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_136  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_137  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_138  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_139  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_140  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_141  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_142  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_143  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_144  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_145  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_146  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_147  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_148  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_149  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_150  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_151  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_152  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_153  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_154  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_155  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_156  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_157  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_158  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_159  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_160  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_161  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_162  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_163  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_164  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_165  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_166  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_167  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_168  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_169  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_170  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_171  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_172  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_173  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_174  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_175  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_176  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_177  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_178  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_179  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_180  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_181  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_182  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_183  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_184  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_185  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_186  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_187  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_188  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_189  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_190  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_191  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_192  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_193  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_194  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_195  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_196  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_197  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_198  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_199  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_200  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_201  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_202  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_203  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_204  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_205  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_206  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_207  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_208  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_209  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_210  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_211  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_212  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_213  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_214  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_215  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_216  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_217  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_218  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_219  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_220  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_221  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_222  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_223  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_224  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_225  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_226  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_227  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_228  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_229  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_230  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_231  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_232  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_233  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_234  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_235  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_236  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_237  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_238  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_239  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_240  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_241  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_242  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_243  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_244  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_245  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_246  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_247  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_248  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_249  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_250  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_251  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_252  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_253  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_254  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_255  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_256  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_257  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_258  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_259  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_260  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_261  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_262  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_263  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_264  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_265  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_266  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_267  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_268  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_269  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_270  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_271  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_272  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_273  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_274  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_275  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_276  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_277  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_278  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_279  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_280  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_281  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_282  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_283  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_284  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_285  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_286  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_287  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_288  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_289  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_290  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_291  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_292  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_293  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_294  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_295  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_296  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_297  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_298  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_299  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_300  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_301  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_302  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_303  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_304  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_305  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_306  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_307  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_308  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_309  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_310  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_311  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_312  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_313  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_314  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_315  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_316  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_317  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_318  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_319  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_320  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_321  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_322  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_323  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_324  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_325  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_326  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_327  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_328  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_329  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_330  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_331  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_332  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_333  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_334  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_335  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_336  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_337  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_338  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_339  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_340  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_341  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_342  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_343  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_344  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_345  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_346  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_347  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_348  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_349  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_350  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_351  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_352  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_353  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_354  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_355  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_356  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_357  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_358  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_359  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_360  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_361  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_362  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_363  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_364  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_365  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_366  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_367  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_368  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_369  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_370  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_371  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_372  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_373  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_374  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_375  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_376  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_377  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_378  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_379  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_380  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_381  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_382  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_383  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_384  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_385  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_386  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_387  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_388  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_389  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_390  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_391  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_392  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_393  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_394  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_395  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_396  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_397  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_398  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_399  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_400  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_401  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_402  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_403  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_404  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_405  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_406  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_407  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_408  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_409  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_410  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_411  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_412  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_413  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_414  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_415  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_416  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_417  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_418  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_419  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_420  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_421  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_422  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_423  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_424  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_425  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_426  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_427  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_428  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_429  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_430  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_431  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_432  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_433  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_434  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_435  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_436  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_437  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_438  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_439  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_440  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_441  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_442  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_443  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_444  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_445  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_446  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_447  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_448  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_449  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_450  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_451  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_452  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_453  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_454  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_455  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_456  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_457  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_458  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_459  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_460  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_461  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_462  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_463  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_464  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_465  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_466  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_467  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_468  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_469  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_470  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_471  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_472  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_473  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_474  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_475  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_476  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_477  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_478  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_479  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_480  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_481  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_482  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_483  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_484  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_485  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_486  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_487  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_488  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_489  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_490  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_491  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_492  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_493  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_494  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_495  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_496  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_497  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_498  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_499  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_500  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_501  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_502  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_503  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_504  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_505  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_506  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_507  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_508  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_509  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_510  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_511  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_512  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_513  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_514  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_515  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_516  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_517  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_518  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_519  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_520  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_521  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_522  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_523  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_524  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_525  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_526  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_527  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_528  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_529  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_530  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_531  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_532  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_533  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_534  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_535  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_536  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_537  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_538  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_539  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_540  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_541  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_542  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_543  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_544  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_545  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_546  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_547  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_548  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_549  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_550  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_551  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_552  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_553  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_554  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_555  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_556  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_557  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_558  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_559  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_560  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_561  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_562  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_563  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_564  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_565  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_566  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_567  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_568  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_569  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_570  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_571  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_572  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_573  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_574  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_575  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_576  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_577  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_578  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_579  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_580  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_581  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_582  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_583  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_584  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_585  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_586  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_587  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_588  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_589  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_590  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_591  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_592  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_593  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_594  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_595  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_596  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_597  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_598  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_599  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_600  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_601  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_602  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_603  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_604  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_605  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_606  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_607  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_608  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_609  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_610  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_611  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_612  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_613  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_614  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_615  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_616  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_617  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_618  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_619  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_620  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_621  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_622  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_623  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_624  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_625  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_626  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_627  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_628  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_629  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_630  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_631  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_632  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_633  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_634  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_635  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_636  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_637  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_638  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_639  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_640  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_641  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_642  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_643  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_644  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_645  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_646  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_647  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_648  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_649  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_650  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_651  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_652  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_653  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_654  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_655  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_656  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_657  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_658  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_659  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_660  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_661  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_662  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_663  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_664  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_665  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_666  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_667  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_668  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_669  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_670  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_671  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_672  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_673  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_674  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_675  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_676  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_677  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_678  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_679  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_680  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_681  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_682  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_683  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_684  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_685  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_686  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_687  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_688  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_689  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_690  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_691  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_692  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_693  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_694  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_695  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_696  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_697  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_698  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_699  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_700  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_701  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_702  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_703  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_704  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_705  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_706  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_707  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_708  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_709  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_710  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_711  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_712  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_713  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_714  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_715  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_716  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_717  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_718  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_719  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_720  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_721  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_722  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_723  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_724  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_725  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_726  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_727  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_728  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_729  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_730  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_731  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_732  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_733  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_734  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_735  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_736  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_737  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_738  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_739  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_740  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_741  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_742  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_743  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_744  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_745  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_746  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_747  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_748  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_749  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_750  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_751  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_752  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_753  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_754  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_755  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_756  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_757  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_758  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_759  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_760  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_761  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_762  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_763  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_764  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_765  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_766  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_767  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_768  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_769  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_770  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_771  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_772  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_773  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_774  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_775  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_776  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_777  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_778  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_779  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_780  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_781  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_782  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_783  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_784  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_785  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_786  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_787  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_788  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_789  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_790  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_791  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_792  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_793  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_794  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_795  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_796  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_797  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_798  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_799  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_800  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_801  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_802  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_803  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_804  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_805  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_806  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_807  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_808  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_809  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_810  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_811  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_812  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_813  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_814  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_815  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_816  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_817  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_818  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_819  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_820  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_821  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_822  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_823  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_824  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_825  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_826  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_827  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_828  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_829  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_830  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_831  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_832  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_833  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_834  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_835  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_836  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_837  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_838  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_839  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_840  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_841  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_842  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_843  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_844  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_845  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_846  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_847  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_848  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_849  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_850  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_851  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_852  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_853  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_854  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_855  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_856  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_857  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_858  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_859  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_860  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_861  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_862  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_863  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_864  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_865  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_866  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_867  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_868  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_869  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_870  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_871  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_872  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_873  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_874  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_875  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_876  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_877  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_878  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_879  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_880  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_881  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_882  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_883  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_884  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_885  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_886  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_887  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_888  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_889  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_890  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_891  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_892  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_893  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_894  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_895  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_896  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_897  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_898  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_899  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_900  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_901  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_902  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_903  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_904  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_905  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_906  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_907  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_908  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_909  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_910  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_911  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_912  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_913  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_914  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_915  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_916  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_917  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_918  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_919  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_920  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_921  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_922  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_923  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_924  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_925  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_926  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_927  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_928  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_929  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_930  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_931  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_932  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_933  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_934  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_935  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_936  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_937  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_938  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_939  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_940  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_941  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_942  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_943  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_944  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_945  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_946  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_947  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_948  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_949  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_950  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_951  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_952  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_953  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_954  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_955  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_956  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_957  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_958  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_959  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_960  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_961  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_962  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_963  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_964  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_965  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_966  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_967  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_968  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_969  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_970  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_971  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_972  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_973  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_974  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_975  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_976  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_977  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_978  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_979  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_980  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_981  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_982  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_983  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_984  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_985  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_986  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_987  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_988  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_989  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_990  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_991  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_992  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_993  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_994  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_995  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_996  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_997  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_998  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_999  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1000 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1001 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1002 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1003 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1004 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1005 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1006 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1007 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1008 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1009 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1010 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1011 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1012 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1013 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1014 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1015 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1016 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1017 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1018 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1019 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1020 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1021 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1022 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1023 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_1024 :out std_logic_vector(11 downto 0);
	   
	   o_Energy_Bin_Pos_1    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_2    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_3    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_4    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_5    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_6    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_7    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_8    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_9    :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_10   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_11   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_12   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_13   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_14   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_15   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_16   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_17   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_18   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_19   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_20   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_21   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_22   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_23   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_24   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_25   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_26   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_27   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_28   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_29   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_30   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_31   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_32   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_33   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_34   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_35   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_36   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_37   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_38   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_39   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_40   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_41   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_42   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_43   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_44   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_45   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_46   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_47   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_48   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_49   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_50   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_51   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_52   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_53   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_54   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_55   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_56   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_57   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_58   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_59   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_60   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_61   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_62   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_63   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_64   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_65   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_66   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_67   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_68   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_69   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_70   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_71   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_72   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_73   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_74   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_75   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_76   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_77   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_78   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_79   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_80   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_81   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_82   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_83   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_84   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_85   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_86   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_87   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_88   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_89   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_90   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_91   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_92   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_93   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_94   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_95   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_96   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_97   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_98   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_99   :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_100  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_101  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_102  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_103  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_104  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_105  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_106  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_107  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_108  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_109  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_110  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_111  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_112  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_113  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_114  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_115  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_116  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_117  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_118  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_119  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_120  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_121  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_122  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_123  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_124  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_125  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_126  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_127  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_128  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_129  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_130  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_131  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_132  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_133  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_134  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_135  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_136  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_137  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_138  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_139  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_140  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_141  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_142  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_143  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_144  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_145  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_146  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_147  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_148  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_149  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_150  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_151  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_152  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_153  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_154  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_155  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_156  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_157  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_158  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_159  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_160  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_161  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_162  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_163  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_164  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_165  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_166  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_167  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_168  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_169  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_170  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_171  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_172  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_173  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_174  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_175  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_176  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_177  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_178  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_179  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_180  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_181  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_182  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_183  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_184  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_185  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_186  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_187  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_188  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_189  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_190  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_191  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_192  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_193  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_194  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_195  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_196  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_197  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_198  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_199  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_200  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_201  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_202  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_203  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_204  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_205  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_206  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_207  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_208  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_209  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_210  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_211  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_212  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_213  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_214  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_215  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_216  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_217  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_218  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_219  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_220  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_221  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_222  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_223  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_224  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_225  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_226  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_227  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_228  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_229  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_230  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_231  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_232  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_233  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_234  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_235  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_236  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_237  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_238  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_239  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_240  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_241  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_242  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_243  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_244  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_245  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_246  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_247  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_248  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_249  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_250  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_251  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_252  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_253  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_254  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_255  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_256  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_257  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_258  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_259  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_260  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_261  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_262  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_263  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_264  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_265  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_266  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_267  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_268  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_269  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_270  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_271  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_272  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_273  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_274  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_275  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_276  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_277  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_278  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_279  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_280  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_281  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_282  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_283  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_284  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_285  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_286  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_287  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_288  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_289  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_290  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_291  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_292  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_293  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_294  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_295  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_296  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_297  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_298  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_299  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_300  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_301  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_302  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_303  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_304  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_305  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_306  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_307  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_308  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_309  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_310  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_311  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_312  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_313  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_314  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_315  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_316  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_317  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_318  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_319  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_320  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_321  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_322  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_323  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_324  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_325  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_326  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_327  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_328  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_329  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_330  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_331  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_332  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_333  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_334  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_335  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_336  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_337  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_338  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_339  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_340  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_341  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_342  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_343  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_344  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_345  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_346  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_347  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_348  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_349  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_350  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_351  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_352  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_353  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_354  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_355  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_356  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_357  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_358  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_359  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_360  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_361  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_362  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_363  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_364  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_365  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_366  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_367  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_368  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_369  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_370  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_371  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_372  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_373  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_374  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_375  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_376  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_377  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_378  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_379  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_380  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_381  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_382  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_383  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_384  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_385  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_386  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_387  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_388  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_389  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_390  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_391  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_392  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_393  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_394  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_395  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_396  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_397  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_398  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_399  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_400  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_401  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_402  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_403  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_404  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_405  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_406  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_407  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_408  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_409  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_410  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_411  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_412  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_413  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_414  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_415  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_416  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_417  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_418  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_419  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_420  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_421  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_422  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_423  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_424  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_425  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_426  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_427  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_428  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_429  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_430  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_431  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_432  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_433  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_434  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_435  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_436  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_437  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_438  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_439  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_440  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_441  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_442  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_443  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_444  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_445  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_446  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_447  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_448  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_449  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_450  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_451  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_452  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_453  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_454  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_455  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_456  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_457  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_458  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_459  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_460  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_461  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_462  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_463  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_464  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_465  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_466  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_467  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_468  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_469  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_470  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_471  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_472  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_473  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_474  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_475  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_476  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_477  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_478  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_479  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_480  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_481  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_482  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_483  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_484  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_485  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_486  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_487  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_488  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_489  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_490  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_491  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_492  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_493  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_494  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_495  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_496  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_497  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_498  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_499  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_500  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_501  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_502  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_503  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_504  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_505  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_506  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_507  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_508  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_509  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_510  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_511  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_512  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_513  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_514  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_515  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_516  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_517  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_518  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_519  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_520  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_521  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_522  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_523  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_524  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_525  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_526  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_527  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_528  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_529  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_530  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_531  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_532  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_533  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_534  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_535  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_536  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_537  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_538  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_539  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_540  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_541  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_542  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_543  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_544  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_545  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_546  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_547  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_548  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_549  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_550  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_551  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_552  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_553  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_554  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_555  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_556  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_557  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_558  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_559  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_560  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_561  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_562  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_563  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_564  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_565  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_566  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_567  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_568  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_569  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_570  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_571  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_572  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_573  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_574  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_575  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_576  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_577  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_578  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_579  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_580  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_581  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_582  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_583  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_584  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_585  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_586  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_587  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_588  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_589  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_590  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_591  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_592  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_593  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_594  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_595  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_596  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_597  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_598  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_599  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_600  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_601  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_602  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_603  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_604  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_605  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_606  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_607  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_608  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_609  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_610  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_611  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_612  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_613  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_614  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_615  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_616  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_617  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_618  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_619  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_620  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_621  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_622  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_623  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_624  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_625  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_626  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_627  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_628  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_629  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_630  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_631  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_632  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_633  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_634  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_635  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_636  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_637  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_638  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_639  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_640  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_641  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_642  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_643  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_644  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_645  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_646  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_647  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_648  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_649  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_650  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_651  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_652  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_653  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_654  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_655  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_656  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_657  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_658  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_659  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_660  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_661  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_662  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_663  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_664  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_665  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_666  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_667  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_668  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_669  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_670  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_671  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_672  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_673  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_674  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_675  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_676  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_677  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_678  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_679  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_680  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_681  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_682  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_683  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_684  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_685  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_686  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_687  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_688  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_689  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_690  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_691  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_692  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_693  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_694  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_695  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_696  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_697  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_698  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_699  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_700  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_701  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_702  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_703  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_704  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_705  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_706  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_707  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_708  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_709  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_710  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_711  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_712  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_713  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_714  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_715  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_716  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_717  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_718  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_719  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_720  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_721  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_722  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_723  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_724  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_725  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_726  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_727  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_728  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_729  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_730  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_731  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_732  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_733  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_734  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_735  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_736  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_737  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_738  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_739  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_740  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_741  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_742  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_743  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_744  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_745  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_746  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_747  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_748  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_749  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_750  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_751  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_752  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_753  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_754  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_755  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_756  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_757  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_758  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_759  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_760  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_761  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_762  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_763  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_764  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_765  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_766  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_767  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_768  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_769  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_770  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_771  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_772  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_773  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_774  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_775  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_776  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_777  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_778  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_779  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_780  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_781  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_782  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_783  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_784  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_785  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_786  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_787  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_788  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_789  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_790  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_791  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_792  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_793  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_794  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_795  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_796  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_797  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_798  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_799  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_800  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_801  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_802  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_803  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_804  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_805  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_806  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_807  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_808  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_809  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_810  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_811  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_812  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_813  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_814  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_815  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_816  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_817  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_818  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_819  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_820  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_821  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_822  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_823  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_824  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_825  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_826  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_827  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_828  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_829  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_830  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_831  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_832  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_833  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_834  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_835  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_836  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_837  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_838  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_839  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_840  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_841  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_842  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_843  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_844  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_845  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_846  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_847  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_848  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_849  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_850  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_851  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_852  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_853  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_854  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_855  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_856  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_857  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_858  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_859  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_860  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_861  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_862  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_863  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_864  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_865  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_866  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_867  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_868  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_869  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_870  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_871  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_872  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_873  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_874  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_875  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_876  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_877  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_878  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_879  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_880  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_881  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_882  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_883  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_884  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_885  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_886  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_887  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_888  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_889  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_890  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_891  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_892  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_893  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_894  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_895  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_896  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_897  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_898  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_899  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_900  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_901  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_902  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_903  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_904  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_905  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_906  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_907  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_908  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_909  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_910  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_911  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_912  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_913  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_914  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_915  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_916  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_917  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_918  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_919  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_920  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_921  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_922  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_923  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_924  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_925  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_926  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_927  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_928  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_929  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_930  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_931  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_932  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_933  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_934  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_935  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_936  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_937  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_938  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_939  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_940  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_941  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_942  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_943  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_944  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_945  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_946  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_947  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_948  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_949  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_950  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_951  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_952  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_953  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_954  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_955  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_956  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_957  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_958  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_959  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_960  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_961  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_962  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_963  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_964  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_965  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_966  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_967  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_968  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_969  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_970  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_971  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_972  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_973  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_974  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_975  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_976  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_977  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_978  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_979  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_980  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_981  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_982  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_983  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_984  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_985  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_986  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_987  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_988  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_989  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_990  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_991  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_992  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_993  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_994  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_995  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_996  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_997  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_998  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_999  :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1000 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1001 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1002 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1003 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1004 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1005 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1006 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1007 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1008 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1009 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1010 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1011 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1012 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1013 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1014 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1015 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1016 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1017 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1018 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1019 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1020 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1021 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1022 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1023 :out std_logic_vector(11 downto 0);
	   o_Energy_Bin_Pos_1024 :out std_logic_vector(11 downto 0)

       );

end entity;
--============================================================================
-- Entity declaration section end
--****************************************************************************


--****************************************************************************
-- Architecture definition section start - RTL
--============================================================================
architecture PeakDetector_RTL of PeakDetector is
attribute syn_preserve : boolean;
attribute syn_preserve of PeakDetector_RTL: architecture is true;

                      
  signal DataRdy_s    :std_logic:='0'; /* synthesis preserve=1*/
  signal DataRdyRis_s :std_logic:='0'; /* synthesis preserve=1*/       

  -- data registers
  signal Data0_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0) 
                          :=(others =>'0'); /* synthesis preserve=1*/
  signal Data1_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/
						  
  signal Data2_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/       
  signal Data3_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data4_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data5_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/                          
  signal Data6_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/    
  signal Data7_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data8_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data9_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/ 
  signal Data10_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/ 
  signal Data11_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/  	
						  
  signal Data12_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/
						  
						  
  signal Data13_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/
  signal Data14_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/       
  signal Data15_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data16_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data17_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/                          
  signal Data18_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/    
  signal Data19_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data20_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data21_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/ 
  signal Data22_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/ 
						  
  signal Data23_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/ 
  signal Data24_s_C1       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/  		
                        				  
						  
  signal Data0_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/
  signal Data1_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/
						  
  signal Data2_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/        
  signal Data3_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data4_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data5_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/                          
  signal Data6_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/    
  signal Data7_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data8_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data9_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/ 
  signal Data10_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data11_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/  	
						  
  signal Data12_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/
						  
						  
  signal Data13_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/
  signal Data14_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/       
  signal Data15_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data16_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data17_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/                          
  signal Data18_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/    
  signal Data19_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data20_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/   
  signal Data21_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/ 
  signal Data22_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/  	
  signal Data23_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/  
  signal Data24_s_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0'); /* synthesis preserve=1*/ 

  signal s_DATA_OUT_C1    :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0');   
  signal s_DATA_OUT_C2       :std_logic_vector(WdVecSize_g-5 downto 0)
                          :=(others =>'0');   
  signal PEAK_C1              :std_logic_vector(11 downto 0)	    :=(others =>'0');
  signal PEAK_C2              :std_logic_vector(11 downto 0)	    :=(others =>'0');	                         				
  signal PEAK_C1_pos          :std_logic_vector(11 downto 0)	    :=(others =>'0');
  signal PEAK_C2_pos          :std_logic_vector(11 downto 0)	    :=(others =>'0');		  

  signal s_PEAK_THD       	  : std_logic_vector(11 downto 0);
  signal s_PEAK_THD_pos       : std_logic_vector(11 downto 0);
  
  signal Energy_Bin_Rdy       :std_logic:='0';
  signal Energy_Bin_Rdy_pos   :std_logic:='0';
  
  signal Energy_Bin_Rdy_bk    :std_logic:='0';
  signal Energy_Bin_Rdy_wr    :std_logic:='0';
  
  
signal s_Energy_Bin_1     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_2     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_3     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_4     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_5     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_6     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_7     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_8     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_9     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_10    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_11    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_12    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_13    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_14    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_15    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_16    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_17    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_18    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_19    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_20    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_21    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_22    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_23    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_24    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_25    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_26    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_27    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_28    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_29    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_30    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_31    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_32    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_33    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_34    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_35    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_36    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_37    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_38    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_39    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_40    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_41    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_42    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_43    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_44    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_45    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_46    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_47    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_48    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_49    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_50    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_51    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_52    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_53    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_54    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_55    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_56    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_57    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_58    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_59    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_60    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_61    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_62    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_63    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_64    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_65    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_66    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_67    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_68    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_69    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_70    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_71    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_72    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_73    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_74    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_75    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_76    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_77    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_78    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_79    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_80    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_81    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_82    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_83    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_84    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_85    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_86    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_87    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_88    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_89    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_90    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_91    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_92    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_93    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_94    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_95    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_96    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_97    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_98    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_99    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_100   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_101   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_102   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_103   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_104   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_105   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_106   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_107   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_108   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_109   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_110   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_111   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_112   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_113   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_114   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_115   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_116   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_117   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_118   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_119   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_120   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_121   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_122   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_123   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_124   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_125   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_126   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_127   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_128   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_129   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_130   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_131   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_132   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_133   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_134   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_135   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_136   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_137   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_138   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_139   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_140   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_141   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_142   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_143   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_144   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_145   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_146   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_147   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_148   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_149   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_150   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_151   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_152   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_153   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_154   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_155   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_156   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_157   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_158   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_159   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_160   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_161   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_162   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_163   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_164   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_165   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_166   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_167   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_168   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_169   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_170   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_171   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_172   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_173   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_174   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_175   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_176   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_177   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_178   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_179   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_180   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_181   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_182   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_183   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_184   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_185   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_186   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_187   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_188   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_189   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_190   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_191   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_192   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_193   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_194   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_195   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_196   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_197   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_198   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_199   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_200   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_201   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_202   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_203   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_204   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_205   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_206   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_207   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_208   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_209   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_210   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_211   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_212   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_213   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_214   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_215   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_216   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_217   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_218   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_219   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_220   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_221   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_222   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_223   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_224   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_225   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_226   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_227   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_228   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_229   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_230   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_231   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_232   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_233   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_234   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_235   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_236   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_237   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_238   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_239   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_240   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_241   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_242   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_243   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_244   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_245   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_246   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_247   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_248   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_249   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_250   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_251   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_252   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_253   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_254   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_255   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_256   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_257   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_258   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_259   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_260   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_261   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_262   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_263   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_264   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_265   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_266   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_267   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_268   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_269   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_270   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_271   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_272   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_273   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_274   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_275   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_276   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_277   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_278   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_279   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_280   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_281   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_282   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_283   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_284   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_285   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_286   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_287   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_288   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_289   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_290   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_291   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_292   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_293   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_294   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_295   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_296   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_297   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_298   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_299   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_300   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_301   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_302   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_303   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_304   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_305   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_306   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_307   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_308   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_309   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_310   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_311   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_312   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_313   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_314   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_315   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_316   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_317   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_318   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_319   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_320   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_321   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_322   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_323   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_324   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_325   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_326   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_327   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_328   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_329   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_330   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_331   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_332   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_333   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_334   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_335   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_336   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_337   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_338   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_339   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_340   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_341   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_342   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_343   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_344   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_345   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_346   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_347   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_348   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_349   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_350   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_351   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_352   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_353   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_354   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_355   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_356   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_357   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_358   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_359   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_360   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_361   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_362   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_363   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_364   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_365   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_366   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_367   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_368   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_369   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_370   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_371   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_372   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_373   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_374   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_375   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_376   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_377   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_378   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_379   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_380   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_381   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_382   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_383   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_384   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_385   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_386   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_387   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_388   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_389   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_390   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_391   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_392   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_393   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_394   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_395   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_396   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_397   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_398   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_399   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_400   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_401   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_402   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_403   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_404   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_405   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_406   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_407   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_408   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_409   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_410   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_411   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_412   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_413   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_414   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_415   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_416   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_417   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_418   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_419   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_420   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_421   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_422   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_423   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_424   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_425   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_426   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_427   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_428   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_429   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_430   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_431   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_432   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_433   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_434   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_435   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_436   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_437   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_438   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_439   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_440   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_441   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_442   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_443   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_444   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_445   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_446   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_447   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_448   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_449   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_450   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_451   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_452   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_453   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_454   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_455   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_456   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_457   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_458   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_459   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_460   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_461   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_462   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_463   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_464   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_465   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_466   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_467   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_468   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_469   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_470   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_471   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_472   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_473   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_474   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_475   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_476   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_477   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_478   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_479   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_480   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_481   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_482   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_483   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_484   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_485   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_486   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_487   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_488   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_489   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_490   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_491   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_492   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_493   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_494   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_495   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_496   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_497   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_498   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_499   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_500   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_501   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_502   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_503   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_504   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_505   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_506   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_507   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_508   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_509   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_510   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_511   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_512   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_513   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_514   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_515   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_516   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_517   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_518   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_519   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_520   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_521   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_522   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_523   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_524   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_525   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_526   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_527   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_528   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_529   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_530   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_531   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_532   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_533   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_534   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_535   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_536   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_537   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_538   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_539   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_540   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_541   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_542   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_543   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_544   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_545   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_546   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_547   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_548   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_549   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_550   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_551   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_552   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_553   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_554   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_555   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_556   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_557   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_558   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_559   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_560   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_561   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_562   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_563   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_564   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_565   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_566   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_567   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_568   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_569   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_570   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_571   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_572   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_573   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_574   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_575   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_576   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_577   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_578   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_579   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_580   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_581   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_582   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_583   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_584   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_585   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_586   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_587   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_588   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_589   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_590   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_591   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_592   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_593   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_594   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_595   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_596   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_597   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_598   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_599   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_600   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_601   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_602   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_603   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_604   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_605   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_606   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_607   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_608   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_609   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_610   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_611   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_612   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_613   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_614   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_615   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_616   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_617   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_618   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_619   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_620   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_621   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_622   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_623   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_624   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_625   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_626   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_627   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_628   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_629   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_630   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_631   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_632   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_633   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_634   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_635   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_636   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_637   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_638   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_639   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_640   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_641   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_642   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_643   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_644   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_645   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_646   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_647   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_648   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_649   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_650   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_651   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_652   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_653   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_654   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_655   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_656   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_657   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_658   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_659   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_660   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_661   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_662   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_663   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_664   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_665   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_666   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_667   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_668   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_669   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_670   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_671   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_672   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_673   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_674   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_675   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_676   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_677   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_678   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_679   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_680   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_681   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_682   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_683   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_684   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_685   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_686   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_687   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_688   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_689   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_690   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_691   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_692   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_693   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_694   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_695   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_696   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_697   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_698   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_699   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_700   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_701   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_702   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_703   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_704   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_705   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_706   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_707   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_708   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_709   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_710   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_711   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_712   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_713   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_714   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_715   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_716   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_717   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_718   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_719   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_720   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_721   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_722   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_723   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_724   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_725   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_726   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_727   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_728   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_729   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_730   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_731   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_732   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_733   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_734   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_735   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_736   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_737   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_738   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_739   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_740   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_741   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_742   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_743   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_744   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_745   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_746   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_747   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_748   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_749   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_750   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_751   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_752   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_753   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_754   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_755   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_756   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_757   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_758   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_759   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_760   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_761   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_762   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_763   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_764   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_765   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_766   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_767   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_768   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_769   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_770   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_771   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_772   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_773   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_774   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_775   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_776   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_777   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_778   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_779   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_780   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_781   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_782   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_783   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_784   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_785   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_786   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_787   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_788   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_789   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_790   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_791   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_792   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_793   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_794   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_795   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_796   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_797   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_798   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_799   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_800   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_801   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_802   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_803   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_804   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_805   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_806   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_807   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_808   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_809   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_810   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_811   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_812   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_813   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_814   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_815   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_816   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_817   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_818   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_819   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_820   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_821   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_822   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_823   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_824   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_825   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_826   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_827   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_828   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_829   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_830   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_831   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_832   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_833   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_834   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_835   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_836   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_837   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_838   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_839   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_840   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_841   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_842   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_843   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_844   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_845   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_846   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_847   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_848   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_849   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_850   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_851   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_852   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_853   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_854   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_855   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_856   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_857   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_858   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_859   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_860   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_861   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_862   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_863   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_864   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_865   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_866   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_867   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_868   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_869   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_870   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_871   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_872   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_873   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_874   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_875   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_876   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_877   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_878   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_879   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_880   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_881   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_882   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_883   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_884   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_885   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_886   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_887   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_888   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_889   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_890   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_891   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_892   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_893   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_894   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_895   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_896   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_897   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_898   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_899   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_900   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_901   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_902   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_903   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_904   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_905   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_906   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_907   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_908   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_909   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_910   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_911   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_912   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_913   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_914   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_915   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_916   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_917   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_918   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_919   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_920   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_921   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_922   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_923   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_924   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_925   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_926   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_927   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_928   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_929   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_930   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_931   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_932   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_933   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_934   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_935   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_936   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_937   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_938   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_939   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_940   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_941   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_942   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_943   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_944   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_945   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_946   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_947   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_948   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_949   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_950   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_951   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_952   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_953   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_954   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_955   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_956   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_957   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_958   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_959   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_960   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_961   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_962   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_963   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_964   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_965   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_966   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_967   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_968   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_969   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_970   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_971   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_972   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_973   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_974   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_975   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_976   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_977   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_978   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_979   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_980   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_981   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_982   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_983   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_984   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_985   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_986   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_987   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_988   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_989   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_990   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_991   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_992   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_993   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_994   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_995   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_996   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_997   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_998   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_999   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1000  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1001  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1002  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1003  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1004  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1005  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1006  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1007  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1008  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1009  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1010  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1011  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1012  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1013  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1014  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1015  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1016  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1017  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1018  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1019  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1020  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1021  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1022  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1023  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_1024  :std_logic_vector(11 downto 0);
  
signal s_Energy_Bin_Pos_1     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_2     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_3     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_4     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_5     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_6     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_7     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_8     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_9     :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_10    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_11    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_12    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_13    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_14    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_15    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_16    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_17    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_18    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_19    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_20    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_21    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_22    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_23    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_24    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_25    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_26    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_27    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_28    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_29    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_30    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_31    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_32    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_33    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_34    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_35    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_36    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_37    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_38    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_39    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_40    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_41    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_42    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_43    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_44    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_45    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_46    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_47    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_48    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_49    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_50    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_51    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_52    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_53    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_54    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_55    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_56    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_57    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_58    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_59    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_60    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_61    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_62    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_63    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_64    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_65    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_66    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_67    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_68    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_69    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_70    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_71    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_72    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_73    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_74    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_75    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_76    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_77    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_78    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_79    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_80    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_81    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_82    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_83    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_84    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_85    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_86    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_87    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_88    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_89    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_90    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_91    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_92    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_93    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_94    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_95    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_96    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_97    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_98    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_99    :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_100   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_101   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_102   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_103   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_104   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_105   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_106   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_107   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_108   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_109   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_110   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_111   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_112   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_113   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_114   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_115   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_116   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_117   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_118   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_119   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_120   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_121   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_122   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_123   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_124   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_125   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_126   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_127   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_128   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_129   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_130   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_131   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_132   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_133   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_134   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_135   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_136   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_137   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_138   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_139   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_140   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_141   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_142   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_143   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_144   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_145   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_146   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_147   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_148   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_149   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_150   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_151   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_152   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_153   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_154   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_155   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_156   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_157   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_158   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_159   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_160   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_161   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_162   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_163   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_164   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_165   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_166   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_167   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_168   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_169   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_170   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_171   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_172   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_173   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_174   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_175   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_176   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_177   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_178   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_179   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_180   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_181   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_182   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_183   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_184   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_185   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_186   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_187   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_188   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_189   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_190   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_191   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_192   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_193   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_194   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_195   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_196   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_197   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_198   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_199   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_200   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_201   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_202   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_203   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_204   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_205   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_206   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_207   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_208   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_209   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_210   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_211   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_212   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_213   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_214   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_215   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_216   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_217   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_218   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_219   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_220   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_221   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_222   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_223   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_224   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_225   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_226   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_227   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_228   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_229   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_230   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_231   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_232   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_233   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_234   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_235   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_236   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_237   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_238   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_239   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_240   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_241   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_242   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_243   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_244   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_245   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_246   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_247   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_248   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_249   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_250   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_251   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_252   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_253   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_254   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_255   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_256   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_257   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_258   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_259   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_260   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_261   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_262   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_263   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_264   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_265   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_266   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_267   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_268   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_269   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_270   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_271   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_272   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_273   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_274   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_275   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_276   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_277   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_278   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_279   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_280   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_281   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_282   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_283   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_284   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_285   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_286   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_287   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_288   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_289   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_290   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_291   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_292   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_293   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_294   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_295   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_296   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_297   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_298   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_299   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_300   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_301   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_302   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_303   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_304   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_305   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_306   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_307   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_308   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_309   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_310   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_311   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_312   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_313   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_314   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_315   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_316   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_317   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_318   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_319   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_320   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_321   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_322   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_323   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_324   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_325   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_326   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_327   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_328   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_329   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_330   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_331   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_332   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_333   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_334   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_335   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_336   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_337   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_338   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_339   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_340   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_341   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_342   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_343   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_344   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_345   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_346   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_347   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_348   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_349   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_350   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_351   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_352   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_353   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_354   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_355   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_356   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_357   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_358   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_359   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_360   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_361   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_362   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_363   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_364   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_365   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_366   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_367   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_368   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_369   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_370   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_371   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_372   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_373   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_374   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_375   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_376   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_377   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_378   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_379   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_380   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_381   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_382   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_383   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_384   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_385   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_386   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_387   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_388   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_389   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_390   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_391   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_392   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_393   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_394   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_395   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_396   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_397   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_398   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_399   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_400   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_401   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_402   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_403   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_404   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_405   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_406   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_407   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_408   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_409   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_410   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_411   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_412   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_413   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_414   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_415   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_416   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_417   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_418   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_419   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_420   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_421   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_422   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_423   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_424   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_425   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_426   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_427   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_428   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_429   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_430   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_431   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_432   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_433   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_434   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_435   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_436   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_437   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_438   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_439   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_440   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_441   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_442   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_443   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_444   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_445   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_446   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_447   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_448   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_449   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_450   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_451   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_452   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_453   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_454   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_455   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_456   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_457   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_458   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_459   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_460   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_461   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_462   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_463   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_464   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_465   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_466   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_467   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_468   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_469   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_470   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_471   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_472   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_473   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_474   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_475   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_476   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_477   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_478   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_479   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_480   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_481   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_482   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_483   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_484   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_485   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_486   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_487   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_488   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_489   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_490   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_491   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_492   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_493   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_494   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_495   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_496   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_497   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_498   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_499   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_500   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_501   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_502   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_503   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_504   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_505   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_506   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_507   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_508   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_509   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_510   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_511   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_512   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_513   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_514   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_515   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_516   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_517   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_518   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_519   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_520   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_521   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_522   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_523   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_524   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_525   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_526   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_527   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_528   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_529   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_530   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_531   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_532   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_533   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_534   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_535   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_536   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_537   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_538   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_539   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_540   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_541   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_542   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_543   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_544   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_545   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_546   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_547   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_548   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_549   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_550   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_551   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_552   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_553   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_554   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_555   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_556   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_557   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_558   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_559   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_560   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_561   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_562   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_563   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_564   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_565   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_566   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_567   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_568   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_569   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_570   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_571   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_572   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_573   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_574   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_575   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_576   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_577   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_578   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_579   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_580   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_581   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_582   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_583   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_584   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_585   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_586   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_587   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_588   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_589   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_590   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_591   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_592   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_593   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_594   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_595   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_596   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_597   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_598   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_599   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_600   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_601   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_602   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_603   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_604   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_605   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_606   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_607   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_608   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_609   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_610   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_611   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_612   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_613   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_614   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_615   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_616   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_617   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_618   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_619   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_620   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_621   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_622   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_623   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_624   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_625   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_626   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_627   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_628   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_629   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_630   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_631   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_632   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_633   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_634   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_635   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_636   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_637   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_638   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_639   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_640   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_641   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_642   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_643   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_644   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_645   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_646   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_647   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_648   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_649   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_650   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_651   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_652   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_653   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_654   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_655   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_656   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_657   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_658   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_659   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_660   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_661   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_662   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_663   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_664   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_665   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_666   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_667   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_668   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_669   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_670   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_671   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_672   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_673   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_674   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_675   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_676   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_677   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_678   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_679   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_680   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_681   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_682   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_683   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_684   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_685   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_686   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_687   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_688   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_689   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_690   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_691   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_692   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_693   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_694   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_695   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_696   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_697   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_698   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_699   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_700   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_701   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_702   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_703   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_704   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_705   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_706   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_707   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_708   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_709   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_710   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_711   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_712   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_713   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_714   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_715   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_716   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_717   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_718   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_719   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_720   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_721   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_722   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_723   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_724   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_725   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_726   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_727   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_728   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_729   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_730   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_731   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_732   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_733   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_734   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_735   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_736   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_737   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_738   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_739   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_740   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_741   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_742   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_743   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_744   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_745   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_746   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_747   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_748   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_749   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_750   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_751   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_752   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_753   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_754   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_755   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_756   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_757   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_758   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_759   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_760   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_761   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_762   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_763   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_764   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_765   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_766   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_767   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_768   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_769   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_770   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_771   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_772   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_773   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_774   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_775   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_776   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_777   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_778   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_779   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_780   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_781   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_782   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_783   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_784   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_785   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_786   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_787   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_788   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_789   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_790   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_791   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_792   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_793   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_794   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_795   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_796   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_797   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_798   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_799   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_800   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_801   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_802   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_803   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_804   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_805   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_806   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_807   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_808   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_809   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_810   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_811   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_812   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_813   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_814   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_815   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_816   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_817   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_818   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_819   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_820   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_821   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_822   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_823   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_824   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_825   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_826   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_827   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_828   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_829   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_830   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_831   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_832   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_833   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_834   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_835   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_836   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_837   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_838   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_839   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_840   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_841   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_842   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_843   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_844   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_845   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_846   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_847   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_848   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_849   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_850   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_851   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_852   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_853   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_854   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_855   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_856   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_857   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_858   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_859   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_860   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_861   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_862   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_863   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_864   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_865   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_866   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_867   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_868   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_869   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_870   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_871   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_872   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_873   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_874   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_875   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_876   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_877   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_878   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_879   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_880   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_881   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_882   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_883   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_884   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_885   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_886   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_887   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_888   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_889   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_890   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_891   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_892   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_893   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_894   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_895   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_896   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_897   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_898   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_899   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_900   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_901   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_902   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_903   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_904   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_905   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_906   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_907   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_908   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_909   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_910   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_911   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_912   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_913   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_914   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_915   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_916   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_917   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_918   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_919   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_920   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_921   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_922   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_923   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_924   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_925   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_926   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_927   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_928   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_929   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_930   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_931   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_932   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_933   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_934   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_935   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_936   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_937   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_938   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_939   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_940   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_941   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_942   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_943   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_944   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_945   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_946   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_947   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_948   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_949   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_950   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_951   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_952   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_953   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_954   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_955   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_956   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_957   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_958   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_959   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_960   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_961   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_962   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_963   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_964   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_965   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_966   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_967   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_968   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_969   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_970   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_971   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_972   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_973   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_974   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_975   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_976   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_977   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_978   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_979   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_980   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_981   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_982   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_983   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_984   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_985   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_986   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_987   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_988   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_989   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_990   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_991   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_992   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_993   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_994   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_995   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_996   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_997   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_998   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_999   :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1000  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1001  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1002  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1003  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1004  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1005  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1006  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1007  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1008  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1009  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1010  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1011  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1012  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1013  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1014  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1015  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1016  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1017  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1018  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1019  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1020  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1021  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1022  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1023  :std_logic_vector(11 downto 0);
signal s_Energy_Bin_Pos_1024  :std_logic_vector(11 downto 0);
  
  
  signal Energy_Bin_Pos_Rdy_1	  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_2     :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_3     :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_4     :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_5     :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_6     :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_7     :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_8     :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_9     :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_10    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_11    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_12    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_13    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_14    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_15    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_16    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_17    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_18    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_19    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_20    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_21    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_22    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_23    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_24    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_25    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_26    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_27    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_28    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_29    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_30    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_31    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_32    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_33    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_34    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_35    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_36    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_37    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_38    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_39    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_40    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_41    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_42    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_43    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_44    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_45    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_46    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_47    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_48    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_49    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_50    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_51    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_52    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_53    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_54    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_55    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_56    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_57    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_58    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_59    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_60    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_61    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_62    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_63    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_64    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_65    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_66    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_67    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_68    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_69    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_70    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_71    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_72    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_73    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_74    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_75    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_76    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_77    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_78    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_79    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_80    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_81    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_82    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_83    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_84    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_85    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_86    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_87    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_88    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_89    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_90    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_91    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_92    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_93    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_94    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_95    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_96    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_97    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_98    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_99    :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_100   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_101   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_102   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_103   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_104   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_105   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_106   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_107   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_108   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_109   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_110   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_111   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_112   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_113   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_114   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_115   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_116   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_117   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_118   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_119   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_120   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_121   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_122   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_123   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_124   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_125   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_126   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_127   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_128   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_129   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_130   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_131   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_132   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_133   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_134   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_135   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_136   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_137   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_138   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_139   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_140   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_141   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_142   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_143   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_144   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_145   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_146   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_147   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_148   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_149   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_150   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_151   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_152   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_153   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_154   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_155   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_156   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_157   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_158   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_159   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_160   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_161   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_162   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_163   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_164   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_165   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_166   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_167   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_168   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_169   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_170   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_171   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_172   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_173   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_174   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_175   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_176   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_177   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_178   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_179   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_180   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_181   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_182   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_183   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_184   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_185   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_186   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_187   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_188   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_189   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_190   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_191   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_192   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_193   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_194   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_195   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_196   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_197   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_198   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_199   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_200   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_201   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_202   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_203   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_204   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_205   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_206   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_207   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_208   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_209   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_210   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_211   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_212   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_213   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_214   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_215   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_216   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_217   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_218   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_219   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_220   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_221   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_222   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_223   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_224   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_225   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_226   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_227   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_228   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_229   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_230   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_231   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_232   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_233   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_234   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_235   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_236   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_237   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_238   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_239   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_240   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_241   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_242   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_243   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_244   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_245   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_246   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_247   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_248   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_249   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_250   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_251   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_252   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_253   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_254   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_255   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_256   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_257   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_258   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_259   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_260   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_261   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_262   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_263   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_264   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_265   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_266   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_267   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_268   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_269   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_270   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_271   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_272   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_273   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_274   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_275   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_276   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_277   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_278   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_279   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_280   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_281   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_282   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_283   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_284   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_285   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_286   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_287   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_288   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_289   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_290   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_291   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_292   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_293   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_294   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_295   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_296   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_297   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_298   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_299   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_300   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_301   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_302   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_303   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_304   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_305   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_306   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_307   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_308   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_309   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_310   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_311   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_312   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_313   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_314   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_315   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_316   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_317   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_318   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_319   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_320   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_321   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_322   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_323   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_324   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_325   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_326   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_327   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_328   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_329   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_330   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_331   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_332   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_333   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_334   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_335   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_336   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_337   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_338   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_339   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_340   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_341   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_342   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_343   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_344   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_345   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_346   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_347   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_348   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_349   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_350   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_351   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_352   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_353   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_354   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_355   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_356   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_357   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_358   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_359   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_360   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_361   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_362   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_363   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_364   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_365   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_366   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_367   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_368   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_369   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_370   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_371   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_372   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_373   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_374   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_375   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_376   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_377   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_378   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_379   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_380   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_381   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_382   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_383   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_384   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_385   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_386   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_387   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_388   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_389   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_390   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_391   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_392   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_393   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_394   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_395   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_396   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_397   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_398   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_399   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_400   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_401   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_402   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_403   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_404   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_405   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_406   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_407   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_408   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_409   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_410   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_411   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_412   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_413   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_414   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_415   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_416   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_417   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_418   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_419   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_420   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_421   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_422   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_423   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_424   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_425   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_426   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_427   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_428   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_429   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_430   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_431   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_432   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_433   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_434   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_435   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_436   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_437   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_438   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_439   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_440   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_441   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_442   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_443   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_444   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_445   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_446   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_447   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_448   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_449   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_450   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_451   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_452   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_453   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_454   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_455   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_456   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_457   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_458   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_459   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_460   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_461   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_462   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_463   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_464   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_465   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_466   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_467   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_468   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_469   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_470   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_471   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_472   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_473   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_474   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_475   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_476   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_477   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_478   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_479   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_480   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_481   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_482   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_483   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_484   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_485   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_486   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_487   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_488   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_489   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_490   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_491   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_492   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_493   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_494   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_495   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_496   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_497   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_498   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_499   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_500   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_501   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_502   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_503   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_504   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_505   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_506   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_507   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_508   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_509   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_510   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_511   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_512   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_513   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_514   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_515   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_516   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_517   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_518   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_519   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_520   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_521   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_522   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_523   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_524   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_525   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_526   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_527   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_528   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_529   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_530   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_531   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_532   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_533   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_534   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_535   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_536   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_537   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_538   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_539   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_540   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_541   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_542   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_543   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_544   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_545   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_546   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_547   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_548   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_549   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_550   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_551   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_552   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_553   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_554   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_555   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_556   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_557   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_558   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_559   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_560   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_561   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_562   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_563   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_564   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_565   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_566   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_567   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_568   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_569   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_570   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_571   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_572   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_573   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_574   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_575   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_576   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_577   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_578   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_579   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_580   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_581   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_582   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_583   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_584   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_585   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_586   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_587   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_588   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_589   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_590   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_591   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_592   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_593   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_594   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_595   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_596   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_597   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_598   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_599   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_600   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_601   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_602   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_603   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_604   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_605   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_606   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_607   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_608   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_609   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_610   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_611   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_612   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_613   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_614   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_615   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_616   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_617   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_618   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_619   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_620   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_621   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_622   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_623   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_624   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_625   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_626   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_627   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_628   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_629   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_630   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_631   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_632   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_633   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_634   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_635   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_636   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_637   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_638   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_639   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_640   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_641   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_642   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_643   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_644   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_645   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_646   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_647   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_648   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_649   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_650   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_651   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_652   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_653   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_654   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_655   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_656   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_657   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_658   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_659   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_660   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_661   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_662   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_663   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_664   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_665   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_666   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_667   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_668   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_669   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_670   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_671   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_672   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_673   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_674   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_675   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_676   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_677   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_678   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_679   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_680   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_681   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_682   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_683   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_684   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_685   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_686   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_687   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_688   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_689   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_690   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_691   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_692   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_693   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_694   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_695   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_696   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_697   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_698   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_699   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_700   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_701   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_702   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_703   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_704   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_705   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_706   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_707   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_708   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_709   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_710   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_711   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_712   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_713   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_714   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_715   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_716   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_717   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_718   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_719   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_720   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_721   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_722   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_723   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_724   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_725   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_726   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_727   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_728   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_729   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_730   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_731   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_732   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_733   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_734   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_735   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_736   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_737   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_738   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_739   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_740   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_741   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_742   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_743   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_744   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_745   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_746   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_747   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_748   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_749   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_750   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_751   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_752   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_753   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_754   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_755   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_756   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_757   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_758   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_759   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_760   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_761   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_762   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_763   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_764   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_765   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_766   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_767   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_768   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_769   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_770   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_771   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_772   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_773   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_774   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_775   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_776   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_777   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_778   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_779   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_780   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_781   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_782   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_783   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_784   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_785   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_786   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_787   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_788   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_789   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_790   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_791   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_792   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_793   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_794   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_795   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_796   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_797   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_798   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_799   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_800   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_801   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_802   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_803   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_804   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_805   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_806   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_807   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_808   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_809   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_810   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_811   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_812   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_813   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_814   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_815   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_816   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_817   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_818   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_819   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_820   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_821   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_822   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_823   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_824   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_825   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_826   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_827   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_828   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_829   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_830   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_831   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_832   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_833   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_834   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_835   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_836   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_837   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_838   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_839   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_840   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_841   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_842   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_843   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_844   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_845   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_846   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_847   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_848   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_849   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_850   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_851   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_852   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_853   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_854   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_855   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_856   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_857   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_858   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_859   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_860   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_861   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_862   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_863   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_864   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_865   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_866   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_867   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_868   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_869   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_870   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_871   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_872   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_873   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_874   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_875   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_876   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_877   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_878   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_879   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_880   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_881   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_882   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_883   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_884   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_885   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_886   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_887   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_888   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_889   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_890   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_891   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_892   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_893   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_894   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_895   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_896   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_897   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_898   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_899   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_900   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_901   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_902   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_903   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_904   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_905   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_906   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_907   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_908   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_909   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_910   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_911   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_912   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_913   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_914   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_915   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_916   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_917   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_918   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_919   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_920   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_921   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_922   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_923   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_924   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_925   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_926   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_927   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_928   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_929   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_930   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_931   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_932   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_933   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_934   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_935   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_936   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_937   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_938   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_939   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_940   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_941   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_942   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_943   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_944   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_945   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_946   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_947   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_948   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_949   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_950   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_951   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_952   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_953   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_954   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_955   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_956   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_957   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_958   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_959   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_960   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_961   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_962   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_963   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_964   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_965   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_966   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_967   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_968   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_969   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_970   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_971   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_972   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_973   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_974   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_975   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_976   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_977   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_978   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_979   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_980   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_981   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_982   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_983   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_984   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_985   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_986   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_987   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_988   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_989   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_990   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_991   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_992   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_993   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_994   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_995   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_996   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_997   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_998   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_999   :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1000  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1001  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1002  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1003  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1004  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1005  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1006  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1007  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1008  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1009  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1010  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1011  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1012  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1013  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1014  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1015  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1016  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1017  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1018  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1019  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1020  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1021  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1022  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1023  :std_logic:='0';
  signal Energy_Bin_Pos_Rdy_1024  :std_logic:='0';
  
  signal Energy_Bin_Rdy_1	  :std_logic:='0';
  signal Energy_Bin_Rdy_2     :std_logic:='0';
  signal Energy_Bin_Rdy_3     :std_logic:='0';
  signal Energy_Bin_Rdy_4     :std_logic:='0';
  signal Energy_Bin_Rdy_5     :std_logic:='0';
  signal Energy_Bin_Rdy_6     :std_logic:='0';
  signal Energy_Bin_Rdy_7     :std_logic:='0';
  signal Energy_Bin_Rdy_8     :std_logic:='0';
  signal Energy_Bin_Rdy_9     :std_logic:='0';
  signal Energy_Bin_Rdy_10    :std_logic:='0';
  signal Energy_Bin_Rdy_11    :std_logic:='0';
  signal Energy_Bin_Rdy_12    :std_logic:='0';
  signal Energy_Bin_Rdy_13    :std_logic:='0';
  signal Energy_Bin_Rdy_14    :std_logic:='0';
  signal Energy_Bin_Rdy_15    :std_logic:='0';
  signal Energy_Bin_Rdy_16    :std_logic:='0';
  signal Energy_Bin_Rdy_17    :std_logic:='0';
  signal Energy_Bin_Rdy_18    :std_logic:='0';
  signal Energy_Bin_Rdy_19    :std_logic:='0';
  signal Energy_Bin_Rdy_20    :std_logic:='0';
  signal Energy_Bin_Rdy_21    :std_logic:='0';
  signal Energy_Bin_Rdy_22    :std_logic:='0';
  signal Energy_Bin_Rdy_23    :std_logic:='0';
  signal Energy_Bin_Rdy_24    :std_logic:='0';
  signal Energy_Bin_Rdy_25    :std_logic:='0';
  signal Energy_Bin_Rdy_26    :std_logic:='0';
  signal Energy_Bin_Rdy_27    :std_logic:='0';
  signal Energy_Bin_Rdy_28    :std_logic:='0';
  signal Energy_Bin_Rdy_29    :std_logic:='0';
  signal Energy_Bin_Rdy_30    :std_logic:='0';
  signal Energy_Bin_Rdy_31    :std_logic:='0';
  signal Energy_Bin_Rdy_32    :std_logic:='0';
  signal Energy_Bin_Rdy_33    :std_logic:='0';
  signal Energy_Bin_Rdy_34    :std_logic:='0';
  signal Energy_Bin_Rdy_35    :std_logic:='0';
  signal Energy_Bin_Rdy_36    :std_logic:='0';
  signal Energy_Bin_Rdy_37    :std_logic:='0';
  signal Energy_Bin_Rdy_38    :std_logic:='0';
  signal Energy_Bin_Rdy_39    :std_logic:='0';
  signal Energy_Bin_Rdy_40    :std_logic:='0';
  signal Energy_Bin_Rdy_41    :std_logic:='0';
  signal Energy_Bin_Rdy_42    :std_logic:='0';
  signal Energy_Bin_Rdy_43    :std_logic:='0';
  signal Energy_Bin_Rdy_44    :std_logic:='0';
  signal Energy_Bin_Rdy_45    :std_logic:='0';
  signal Energy_Bin_Rdy_46    :std_logic:='0';
  signal Energy_Bin_Rdy_47    :std_logic:='0';
  signal Energy_Bin_Rdy_48    :std_logic:='0';
  signal Energy_Bin_Rdy_49    :std_logic:='0';
  signal Energy_Bin_Rdy_50    :std_logic:='0';
  signal Energy_Bin_Rdy_51    :std_logic:='0';
  signal Energy_Bin_Rdy_52    :std_logic:='0';
  signal Energy_Bin_Rdy_53    :std_logic:='0';
  signal Energy_Bin_Rdy_54    :std_logic:='0';
  signal Energy_Bin_Rdy_55    :std_logic:='0';
  signal Energy_Bin_Rdy_56    :std_logic:='0';
  signal Energy_Bin_Rdy_57    :std_logic:='0';
  signal Energy_Bin_Rdy_58    :std_logic:='0';
  signal Energy_Bin_Rdy_59    :std_logic:='0';
  signal Energy_Bin_Rdy_60    :std_logic:='0';
  signal Energy_Bin_Rdy_61    :std_logic:='0';
  signal Energy_Bin_Rdy_62    :std_logic:='0';
  signal Energy_Bin_Rdy_63    :std_logic:='0';
  signal Energy_Bin_Rdy_64    :std_logic:='0';
  signal Energy_Bin_Rdy_65    :std_logic:='0';
  signal Energy_Bin_Rdy_66    :std_logic:='0';
  signal Energy_Bin_Rdy_67    :std_logic:='0';
  signal Energy_Bin_Rdy_68    :std_logic:='0';
  signal Energy_Bin_Rdy_69    :std_logic:='0';
  signal Energy_Bin_Rdy_70    :std_logic:='0';
  signal Energy_Bin_Rdy_71    :std_logic:='0';
  signal Energy_Bin_Rdy_72    :std_logic:='0';
  signal Energy_Bin_Rdy_73    :std_logic:='0';
  signal Energy_Bin_Rdy_74    :std_logic:='0';
  signal Energy_Bin_Rdy_75    :std_logic:='0';
  signal Energy_Bin_Rdy_76    :std_logic:='0';
  signal Energy_Bin_Rdy_77    :std_logic:='0';
  signal Energy_Bin_Rdy_78    :std_logic:='0';
  signal Energy_Bin_Rdy_79    :std_logic:='0';
  signal Energy_Bin_Rdy_80    :std_logic:='0';
  signal Energy_Bin_Rdy_81    :std_logic:='0';
  signal Energy_Bin_Rdy_82    :std_logic:='0';
  signal Energy_Bin_Rdy_83    :std_logic:='0';
  signal Energy_Bin_Rdy_84    :std_logic:='0';
  signal Energy_Bin_Rdy_85    :std_logic:='0';
  signal Energy_Bin_Rdy_86    :std_logic:='0';
  signal Energy_Bin_Rdy_87    :std_logic:='0';
  signal Energy_Bin_Rdy_88    :std_logic:='0';
  signal Energy_Bin_Rdy_89    :std_logic:='0';
  signal Energy_Bin_Rdy_90    :std_logic:='0';
  signal Energy_Bin_Rdy_91    :std_logic:='0';
  signal Energy_Bin_Rdy_92    :std_logic:='0';
  signal Energy_Bin_Rdy_93    :std_logic:='0';
  signal Energy_Bin_Rdy_94    :std_logic:='0';
  signal Energy_Bin_Rdy_95    :std_logic:='0';
  signal Energy_Bin_Rdy_96    :std_logic:='0';
  signal Energy_Bin_Rdy_97    :std_logic:='0';
  signal Energy_Bin_Rdy_98    :std_logic:='0';
  signal Energy_Bin_Rdy_99    :std_logic:='0';
  signal Energy_Bin_Rdy_100   :std_logic:='0';
  signal Energy_Bin_Rdy_101   :std_logic:='0';
  signal Energy_Bin_Rdy_102   :std_logic:='0';
  signal Energy_Bin_Rdy_103   :std_logic:='0';
  signal Energy_Bin_Rdy_104   :std_logic:='0';
  signal Energy_Bin_Rdy_105   :std_logic:='0';
  signal Energy_Bin_Rdy_106   :std_logic:='0';
  signal Energy_Bin_Rdy_107   :std_logic:='0';
  signal Energy_Bin_Rdy_108   :std_logic:='0';
  signal Energy_Bin_Rdy_109   :std_logic:='0';
  signal Energy_Bin_Rdy_110   :std_logic:='0';
  signal Energy_Bin_Rdy_111   :std_logic:='0';
  signal Energy_Bin_Rdy_112   :std_logic:='0';
  signal Energy_Bin_Rdy_113   :std_logic:='0';
  signal Energy_Bin_Rdy_114   :std_logic:='0';
  signal Energy_Bin_Rdy_115   :std_logic:='0';
  signal Energy_Bin_Rdy_116   :std_logic:='0';
  signal Energy_Bin_Rdy_117   :std_logic:='0';
  signal Energy_Bin_Rdy_118   :std_logic:='0';
  signal Energy_Bin_Rdy_119   :std_logic:='0';
  signal Energy_Bin_Rdy_120   :std_logic:='0';
  signal Energy_Bin_Rdy_121   :std_logic:='0';
  signal Energy_Bin_Rdy_122   :std_logic:='0';
  signal Energy_Bin_Rdy_123   :std_logic:='0';
  signal Energy_Bin_Rdy_124   :std_logic:='0';
  signal Energy_Bin_Rdy_125   :std_logic:='0';
  signal Energy_Bin_Rdy_126   :std_logic:='0';
  signal Energy_Bin_Rdy_127   :std_logic:='0';
  signal Energy_Bin_Rdy_128   :std_logic:='0';
  signal Energy_Bin_Rdy_129   :std_logic:='0';
  signal Energy_Bin_Rdy_130   :std_logic:='0';
  signal Energy_Bin_Rdy_131   :std_logic:='0';
  signal Energy_Bin_Rdy_132   :std_logic:='0';
  signal Energy_Bin_Rdy_133   :std_logic:='0';
  signal Energy_Bin_Rdy_134   :std_logic:='0';
  signal Energy_Bin_Rdy_135   :std_logic:='0';
  signal Energy_Bin_Rdy_136   :std_logic:='0';
  signal Energy_Bin_Rdy_137   :std_logic:='0';
  signal Energy_Bin_Rdy_138   :std_logic:='0';
  signal Energy_Bin_Rdy_139   :std_logic:='0';
  signal Energy_Bin_Rdy_140   :std_logic:='0';
  signal Energy_Bin_Rdy_141   :std_logic:='0';
  signal Energy_Bin_Rdy_142   :std_logic:='0';
  signal Energy_Bin_Rdy_143   :std_logic:='0';
  signal Energy_Bin_Rdy_144   :std_logic:='0';
  signal Energy_Bin_Rdy_145   :std_logic:='0';
  signal Energy_Bin_Rdy_146   :std_logic:='0';
  signal Energy_Bin_Rdy_147   :std_logic:='0';
  signal Energy_Bin_Rdy_148   :std_logic:='0';
  signal Energy_Bin_Rdy_149   :std_logic:='0';
  signal Energy_Bin_Rdy_150   :std_logic:='0';
  signal Energy_Bin_Rdy_151   :std_logic:='0';
  signal Energy_Bin_Rdy_152   :std_logic:='0';
  signal Energy_Bin_Rdy_153   :std_logic:='0';
  signal Energy_Bin_Rdy_154   :std_logic:='0';
  signal Energy_Bin_Rdy_155   :std_logic:='0';
  signal Energy_Bin_Rdy_156   :std_logic:='0';
  signal Energy_Bin_Rdy_157   :std_logic:='0';
  signal Energy_Bin_Rdy_158   :std_logic:='0';
  signal Energy_Bin_Rdy_159   :std_logic:='0';
  signal Energy_Bin_Rdy_160   :std_logic:='0';
  signal Energy_Bin_Rdy_161   :std_logic:='0';
  signal Energy_Bin_Rdy_162   :std_logic:='0';
  signal Energy_Bin_Rdy_163   :std_logic:='0';
  signal Energy_Bin_Rdy_164   :std_logic:='0';
  signal Energy_Bin_Rdy_165   :std_logic:='0';
  signal Energy_Bin_Rdy_166   :std_logic:='0';
  signal Energy_Bin_Rdy_167   :std_logic:='0';
  signal Energy_Bin_Rdy_168   :std_logic:='0';
  signal Energy_Bin_Rdy_169   :std_logic:='0';
  signal Energy_Bin_Rdy_170   :std_logic:='0';
  signal Energy_Bin_Rdy_171   :std_logic:='0';
  signal Energy_Bin_Rdy_172   :std_logic:='0';
  signal Energy_Bin_Rdy_173   :std_logic:='0';
  signal Energy_Bin_Rdy_174   :std_logic:='0';
  signal Energy_Bin_Rdy_175   :std_logic:='0';
  signal Energy_Bin_Rdy_176   :std_logic:='0';
  signal Energy_Bin_Rdy_177   :std_logic:='0';
  signal Energy_Bin_Rdy_178   :std_logic:='0';
  signal Energy_Bin_Rdy_179   :std_logic:='0';
  signal Energy_Bin_Rdy_180   :std_logic:='0';
  signal Energy_Bin_Rdy_181   :std_logic:='0';
  signal Energy_Bin_Rdy_182   :std_logic:='0';
  signal Energy_Bin_Rdy_183   :std_logic:='0';
  signal Energy_Bin_Rdy_184   :std_logic:='0';
  signal Energy_Bin_Rdy_185   :std_logic:='0';
  signal Energy_Bin_Rdy_186   :std_logic:='0';
  signal Energy_Bin_Rdy_187   :std_logic:='0';
  signal Energy_Bin_Rdy_188   :std_logic:='0';
  signal Energy_Bin_Rdy_189   :std_logic:='0';
  signal Energy_Bin_Rdy_190   :std_logic:='0';
  signal Energy_Bin_Rdy_191   :std_logic:='0';
  signal Energy_Bin_Rdy_192   :std_logic:='0';
  signal Energy_Bin_Rdy_193   :std_logic:='0';
  signal Energy_Bin_Rdy_194   :std_logic:='0';
  signal Energy_Bin_Rdy_195   :std_logic:='0';
  signal Energy_Bin_Rdy_196   :std_logic:='0';
  signal Energy_Bin_Rdy_197   :std_logic:='0';
  signal Energy_Bin_Rdy_198   :std_logic:='0';
  signal Energy_Bin_Rdy_199   :std_logic:='0';
  signal Energy_Bin_Rdy_200   :std_logic:='0';
  signal Energy_Bin_Rdy_201   :std_logic:='0';
  signal Energy_Bin_Rdy_202   :std_logic:='0';
  signal Energy_Bin_Rdy_203   :std_logic:='0';
  signal Energy_Bin_Rdy_204   :std_logic:='0';
  signal Energy_Bin_Rdy_205   :std_logic:='0';
  signal Energy_Bin_Rdy_206   :std_logic:='0';
  signal Energy_Bin_Rdy_207   :std_logic:='0';
  signal Energy_Bin_Rdy_208   :std_logic:='0';
  signal Energy_Bin_Rdy_209   :std_logic:='0';
  signal Energy_Bin_Rdy_210   :std_logic:='0';
  signal Energy_Bin_Rdy_211   :std_logic:='0';
  signal Energy_Bin_Rdy_212   :std_logic:='0';
  signal Energy_Bin_Rdy_213   :std_logic:='0';
  signal Energy_Bin_Rdy_214   :std_logic:='0';
  signal Energy_Bin_Rdy_215   :std_logic:='0';
  signal Energy_Bin_Rdy_216   :std_logic:='0';
  signal Energy_Bin_Rdy_217   :std_logic:='0';
  signal Energy_Bin_Rdy_218   :std_logic:='0';
  signal Energy_Bin_Rdy_219   :std_logic:='0';
  signal Energy_Bin_Rdy_220   :std_logic:='0';
  signal Energy_Bin_Rdy_221   :std_logic:='0';
  signal Energy_Bin_Rdy_222   :std_logic:='0';
  signal Energy_Bin_Rdy_223   :std_logic:='0';
  signal Energy_Bin_Rdy_224   :std_logic:='0';
  signal Energy_Bin_Rdy_225   :std_logic:='0';
  signal Energy_Bin_Rdy_226   :std_logic:='0';
  signal Energy_Bin_Rdy_227   :std_logic:='0';
  signal Energy_Bin_Rdy_228   :std_logic:='0';
  signal Energy_Bin_Rdy_229   :std_logic:='0';
  signal Energy_Bin_Rdy_230   :std_logic:='0';
  signal Energy_Bin_Rdy_231   :std_logic:='0';
  signal Energy_Bin_Rdy_232   :std_logic:='0';
  signal Energy_Bin_Rdy_233   :std_logic:='0';
  signal Energy_Bin_Rdy_234   :std_logic:='0';
  signal Energy_Bin_Rdy_235   :std_logic:='0';
  signal Energy_Bin_Rdy_236   :std_logic:='0';
  signal Energy_Bin_Rdy_237   :std_logic:='0';
  signal Energy_Bin_Rdy_238   :std_logic:='0';
  signal Energy_Bin_Rdy_239   :std_logic:='0';
  signal Energy_Bin_Rdy_240   :std_logic:='0';
  signal Energy_Bin_Rdy_241   :std_logic:='0';
  signal Energy_Bin_Rdy_242   :std_logic:='0';
  signal Energy_Bin_Rdy_243   :std_logic:='0';
  signal Energy_Bin_Rdy_244   :std_logic:='0';
  signal Energy_Bin_Rdy_245   :std_logic:='0';
  signal Energy_Bin_Rdy_246   :std_logic:='0';
  signal Energy_Bin_Rdy_247   :std_logic:='0';
  signal Energy_Bin_Rdy_248   :std_logic:='0';
  signal Energy_Bin_Rdy_249   :std_logic:='0';
  signal Energy_Bin_Rdy_250   :std_logic:='0';
  signal Energy_Bin_Rdy_251   :std_logic:='0';
  signal Energy_Bin_Rdy_252   :std_logic:='0';
  signal Energy_Bin_Rdy_253   :std_logic:='0';
  signal Energy_Bin_Rdy_254   :std_logic:='0';
  signal Energy_Bin_Rdy_255   :std_logic:='0';
  signal Energy_Bin_Rdy_256   :std_logic:='0';
  signal Energy_Bin_Rdy_257   :std_logic:='0';
  signal Energy_Bin_Rdy_258   :std_logic:='0';
  signal Energy_Bin_Rdy_259   :std_logic:='0';
  signal Energy_Bin_Rdy_260   :std_logic:='0';
  signal Energy_Bin_Rdy_261   :std_logic:='0';
  signal Energy_Bin_Rdy_262   :std_logic:='0';
  signal Energy_Bin_Rdy_263   :std_logic:='0';
  signal Energy_Bin_Rdy_264   :std_logic:='0';
  signal Energy_Bin_Rdy_265   :std_logic:='0';
  signal Energy_Bin_Rdy_266   :std_logic:='0';
  signal Energy_Bin_Rdy_267   :std_logic:='0';
  signal Energy_Bin_Rdy_268   :std_logic:='0';
  signal Energy_Bin_Rdy_269   :std_logic:='0';
  signal Energy_Bin_Rdy_270   :std_logic:='0';
  signal Energy_Bin_Rdy_271   :std_logic:='0';
  signal Energy_Bin_Rdy_272   :std_logic:='0';
  signal Energy_Bin_Rdy_273   :std_logic:='0';
  signal Energy_Bin_Rdy_274   :std_logic:='0';
  signal Energy_Bin_Rdy_275   :std_logic:='0';
  signal Energy_Bin_Rdy_276   :std_logic:='0';
  signal Energy_Bin_Rdy_277   :std_logic:='0';
  signal Energy_Bin_Rdy_278   :std_logic:='0';
  signal Energy_Bin_Rdy_279   :std_logic:='0';
  signal Energy_Bin_Rdy_280   :std_logic:='0';
  signal Energy_Bin_Rdy_281   :std_logic:='0';
  signal Energy_Bin_Rdy_282   :std_logic:='0';
  signal Energy_Bin_Rdy_283   :std_logic:='0';
  signal Energy_Bin_Rdy_284   :std_logic:='0';
  signal Energy_Bin_Rdy_285   :std_logic:='0';
  signal Energy_Bin_Rdy_286   :std_logic:='0';
  signal Energy_Bin_Rdy_287   :std_logic:='0';
  signal Energy_Bin_Rdy_288   :std_logic:='0';
  signal Energy_Bin_Rdy_289   :std_logic:='0';
  signal Energy_Bin_Rdy_290   :std_logic:='0';
  signal Energy_Bin_Rdy_291   :std_logic:='0';
  signal Energy_Bin_Rdy_292   :std_logic:='0';
  signal Energy_Bin_Rdy_293   :std_logic:='0';
  signal Energy_Bin_Rdy_294   :std_logic:='0';
  signal Energy_Bin_Rdy_295   :std_logic:='0';
  signal Energy_Bin_Rdy_296   :std_logic:='0';
  signal Energy_Bin_Rdy_297   :std_logic:='0';
  signal Energy_Bin_Rdy_298   :std_logic:='0';
  signal Energy_Bin_Rdy_299   :std_logic:='0';
  signal Energy_Bin_Rdy_300   :std_logic:='0';
  signal Energy_Bin_Rdy_301   :std_logic:='0';
  signal Energy_Bin_Rdy_302   :std_logic:='0';
  signal Energy_Bin_Rdy_303   :std_logic:='0';
  signal Energy_Bin_Rdy_304   :std_logic:='0';
  signal Energy_Bin_Rdy_305   :std_logic:='0';
  signal Energy_Bin_Rdy_306   :std_logic:='0';
  signal Energy_Bin_Rdy_307   :std_logic:='0';
  signal Energy_Bin_Rdy_308   :std_logic:='0';
  signal Energy_Bin_Rdy_309   :std_logic:='0';
  signal Energy_Bin_Rdy_310   :std_logic:='0';
  signal Energy_Bin_Rdy_311   :std_logic:='0';
  signal Energy_Bin_Rdy_312   :std_logic:='0';
  signal Energy_Bin_Rdy_313   :std_logic:='0';
  signal Energy_Bin_Rdy_314   :std_logic:='0';
  signal Energy_Bin_Rdy_315   :std_logic:='0';
  signal Energy_Bin_Rdy_316   :std_logic:='0';
  signal Energy_Bin_Rdy_317   :std_logic:='0';
  signal Energy_Bin_Rdy_318   :std_logic:='0';
  signal Energy_Bin_Rdy_319   :std_logic:='0';
  signal Energy_Bin_Rdy_320   :std_logic:='0';
  signal Energy_Bin_Rdy_321   :std_logic:='0';
  signal Energy_Bin_Rdy_322   :std_logic:='0';
  signal Energy_Bin_Rdy_323   :std_logic:='0';
  signal Energy_Bin_Rdy_324   :std_logic:='0';
  signal Energy_Bin_Rdy_325   :std_logic:='0';
  signal Energy_Bin_Rdy_326   :std_logic:='0';
  signal Energy_Bin_Rdy_327   :std_logic:='0';
  signal Energy_Bin_Rdy_328   :std_logic:='0';
  signal Energy_Bin_Rdy_329   :std_logic:='0';
  signal Energy_Bin_Rdy_330   :std_logic:='0';
  signal Energy_Bin_Rdy_331   :std_logic:='0';
  signal Energy_Bin_Rdy_332   :std_logic:='0';
  signal Energy_Bin_Rdy_333   :std_logic:='0';
  signal Energy_Bin_Rdy_334   :std_logic:='0';
  signal Energy_Bin_Rdy_335   :std_logic:='0';
  signal Energy_Bin_Rdy_336   :std_logic:='0';
  signal Energy_Bin_Rdy_337   :std_logic:='0';
  signal Energy_Bin_Rdy_338   :std_logic:='0';
  signal Energy_Bin_Rdy_339   :std_logic:='0';
  signal Energy_Bin_Rdy_340   :std_logic:='0';
  signal Energy_Bin_Rdy_341   :std_logic:='0';
  signal Energy_Bin_Rdy_342   :std_logic:='0';
  signal Energy_Bin_Rdy_343   :std_logic:='0';
  signal Energy_Bin_Rdy_344   :std_logic:='0';
  signal Energy_Bin_Rdy_345   :std_logic:='0';
  signal Energy_Bin_Rdy_346   :std_logic:='0';
  signal Energy_Bin_Rdy_347   :std_logic:='0';
  signal Energy_Bin_Rdy_348   :std_logic:='0';
  signal Energy_Bin_Rdy_349   :std_logic:='0';
  signal Energy_Bin_Rdy_350   :std_logic:='0';
  signal Energy_Bin_Rdy_351   :std_logic:='0';
  signal Energy_Bin_Rdy_352   :std_logic:='0';
  signal Energy_Bin_Rdy_353   :std_logic:='0';
  signal Energy_Bin_Rdy_354   :std_logic:='0';
  signal Energy_Bin_Rdy_355   :std_logic:='0';
  signal Energy_Bin_Rdy_356   :std_logic:='0';
  signal Energy_Bin_Rdy_357   :std_logic:='0';
  signal Energy_Bin_Rdy_358   :std_logic:='0';
  signal Energy_Bin_Rdy_359   :std_logic:='0';
  signal Energy_Bin_Rdy_360   :std_logic:='0';
  signal Energy_Bin_Rdy_361   :std_logic:='0';
  signal Energy_Bin_Rdy_362   :std_logic:='0';
  signal Energy_Bin_Rdy_363   :std_logic:='0';
  signal Energy_Bin_Rdy_364   :std_logic:='0';
  signal Energy_Bin_Rdy_365   :std_logic:='0';
  signal Energy_Bin_Rdy_366   :std_logic:='0';
  signal Energy_Bin_Rdy_367   :std_logic:='0';
  signal Energy_Bin_Rdy_368   :std_logic:='0';
  signal Energy_Bin_Rdy_369   :std_logic:='0';
  signal Energy_Bin_Rdy_370   :std_logic:='0';
  signal Energy_Bin_Rdy_371   :std_logic:='0';
  signal Energy_Bin_Rdy_372   :std_logic:='0';
  signal Energy_Bin_Rdy_373   :std_logic:='0';
  signal Energy_Bin_Rdy_374   :std_logic:='0';
  signal Energy_Bin_Rdy_375   :std_logic:='0';
  signal Energy_Bin_Rdy_376   :std_logic:='0';
  signal Energy_Bin_Rdy_377   :std_logic:='0';
  signal Energy_Bin_Rdy_378   :std_logic:='0';
  signal Energy_Bin_Rdy_379   :std_logic:='0';
  signal Energy_Bin_Rdy_380   :std_logic:='0';
  signal Energy_Bin_Rdy_381   :std_logic:='0';
  signal Energy_Bin_Rdy_382   :std_logic:='0';
  signal Energy_Bin_Rdy_383   :std_logic:='0';
  signal Energy_Bin_Rdy_384   :std_logic:='0';
  signal Energy_Bin_Rdy_385   :std_logic:='0';
  signal Energy_Bin_Rdy_386   :std_logic:='0';
  signal Energy_Bin_Rdy_387   :std_logic:='0';
  signal Energy_Bin_Rdy_388   :std_logic:='0';
  signal Energy_Bin_Rdy_389   :std_logic:='0';
  signal Energy_Bin_Rdy_390   :std_logic:='0';
  signal Energy_Bin_Rdy_391   :std_logic:='0';
  signal Energy_Bin_Rdy_392   :std_logic:='0';
  signal Energy_Bin_Rdy_393   :std_logic:='0';
  signal Energy_Bin_Rdy_394   :std_logic:='0';
  signal Energy_Bin_Rdy_395   :std_logic:='0';
  signal Energy_Bin_Rdy_396   :std_logic:='0';
  signal Energy_Bin_Rdy_397   :std_logic:='0';
  signal Energy_Bin_Rdy_398   :std_logic:='0';
  signal Energy_Bin_Rdy_399   :std_logic:='0';
  signal Energy_Bin_Rdy_400   :std_logic:='0';
  signal Energy_Bin_Rdy_401   :std_logic:='0';
  signal Energy_Bin_Rdy_402   :std_logic:='0';
  signal Energy_Bin_Rdy_403   :std_logic:='0';
  signal Energy_Bin_Rdy_404   :std_logic:='0';
  signal Energy_Bin_Rdy_405   :std_logic:='0';
  signal Energy_Bin_Rdy_406   :std_logic:='0';
  signal Energy_Bin_Rdy_407   :std_logic:='0';
  signal Energy_Bin_Rdy_408   :std_logic:='0';
  signal Energy_Bin_Rdy_409   :std_logic:='0';
  signal Energy_Bin_Rdy_410   :std_logic:='0';
  signal Energy_Bin_Rdy_411   :std_logic:='0';
  signal Energy_Bin_Rdy_412   :std_logic:='0';
  signal Energy_Bin_Rdy_413   :std_logic:='0';
  signal Energy_Bin_Rdy_414   :std_logic:='0';
  signal Energy_Bin_Rdy_415   :std_logic:='0';
  signal Energy_Bin_Rdy_416   :std_logic:='0';
  signal Energy_Bin_Rdy_417   :std_logic:='0';
  signal Energy_Bin_Rdy_418   :std_logic:='0';
  signal Energy_Bin_Rdy_419   :std_logic:='0';
  signal Energy_Bin_Rdy_420   :std_logic:='0';
  signal Energy_Bin_Rdy_421   :std_logic:='0';
  signal Energy_Bin_Rdy_422   :std_logic:='0';
  signal Energy_Bin_Rdy_423   :std_logic:='0';
  signal Energy_Bin_Rdy_424   :std_logic:='0';
  signal Energy_Bin_Rdy_425   :std_logic:='0';
  signal Energy_Bin_Rdy_426   :std_logic:='0';
  signal Energy_Bin_Rdy_427   :std_logic:='0';
  signal Energy_Bin_Rdy_428   :std_logic:='0';
  signal Energy_Bin_Rdy_429   :std_logic:='0';
  signal Energy_Bin_Rdy_430   :std_logic:='0';
  signal Energy_Bin_Rdy_431   :std_logic:='0';
  signal Energy_Bin_Rdy_432   :std_logic:='0';
  signal Energy_Bin_Rdy_433   :std_logic:='0';
  signal Energy_Bin_Rdy_434   :std_logic:='0';
  signal Energy_Bin_Rdy_435   :std_logic:='0';
  signal Energy_Bin_Rdy_436   :std_logic:='0';
  signal Energy_Bin_Rdy_437   :std_logic:='0';
  signal Energy_Bin_Rdy_438   :std_logic:='0';
  signal Energy_Bin_Rdy_439   :std_logic:='0';
  signal Energy_Bin_Rdy_440   :std_logic:='0';
  signal Energy_Bin_Rdy_441   :std_logic:='0';
  signal Energy_Bin_Rdy_442   :std_logic:='0';
  signal Energy_Bin_Rdy_443   :std_logic:='0';
  signal Energy_Bin_Rdy_444   :std_logic:='0';
  signal Energy_Bin_Rdy_445   :std_logic:='0';
  signal Energy_Bin_Rdy_446   :std_logic:='0';
  signal Energy_Bin_Rdy_447   :std_logic:='0';
  signal Energy_Bin_Rdy_448   :std_logic:='0';
  signal Energy_Bin_Rdy_449   :std_logic:='0';
  signal Energy_Bin_Rdy_450   :std_logic:='0';
  signal Energy_Bin_Rdy_451   :std_logic:='0';
  signal Energy_Bin_Rdy_452   :std_logic:='0';
  signal Energy_Bin_Rdy_453   :std_logic:='0';
  signal Energy_Bin_Rdy_454   :std_logic:='0';
  signal Energy_Bin_Rdy_455   :std_logic:='0';
  signal Energy_Bin_Rdy_456   :std_logic:='0';
  signal Energy_Bin_Rdy_457   :std_logic:='0';
  signal Energy_Bin_Rdy_458   :std_logic:='0';
  signal Energy_Bin_Rdy_459   :std_logic:='0';
  signal Energy_Bin_Rdy_460   :std_logic:='0';
  signal Energy_Bin_Rdy_461   :std_logic:='0';
  signal Energy_Bin_Rdy_462   :std_logic:='0';
  signal Energy_Bin_Rdy_463   :std_logic:='0';
  signal Energy_Bin_Rdy_464   :std_logic:='0';
  signal Energy_Bin_Rdy_465   :std_logic:='0';
  signal Energy_Bin_Rdy_466   :std_logic:='0';
  signal Energy_Bin_Rdy_467   :std_logic:='0';
  signal Energy_Bin_Rdy_468   :std_logic:='0';
  signal Energy_Bin_Rdy_469   :std_logic:='0';
  signal Energy_Bin_Rdy_470   :std_logic:='0';
  signal Energy_Bin_Rdy_471   :std_logic:='0';
  signal Energy_Bin_Rdy_472   :std_logic:='0';
  signal Energy_Bin_Rdy_473   :std_logic:='0';
  signal Energy_Bin_Rdy_474   :std_logic:='0';
  signal Energy_Bin_Rdy_475   :std_logic:='0';
  signal Energy_Bin_Rdy_476   :std_logic:='0';
  signal Energy_Bin_Rdy_477   :std_logic:='0';
  signal Energy_Bin_Rdy_478   :std_logic:='0';
  signal Energy_Bin_Rdy_479   :std_logic:='0';
  signal Energy_Bin_Rdy_480   :std_logic:='0';
  signal Energy_Bin_Rdy_481   :std_logic:='0';
  signal Energy_Bin_Rdy_482   :std_logic:='0';
  signal Energy_Bin_Rdy_483   :std_logic:='0';
  signal Energy_Bin_Rdy_484   :std_logic:='0';
  signal Energy_Bin_Rdy_485   :std_logic:='0';
  signal Energy_Bin_Rdy_486   :std_logic:='0';
  signal Energy_Bin_Rdy_487   :std_logic:='0';
  signal Energy_Bin_Rdy_488   :std_logic:='0';
  signal Energy_Bin_Rdy_489   :std_logic:='0';
  signal Energy_Bin_Rdy_490   :std_logic:='0';
  signal Energy_Bin_Rdy_491   :std_logic:='0';
  signal Energy_Bin_Rdy_492   :std_logic:='0';
  signal Energy_Bin_Rdy_493   :std_logic:='0';
  signal Energy_Bin_Rdy_494   :std_logic:='0';
  signal Energy_Bin_Rdy_495   :std_logic:='0';
  signal Energy_Bin_Rdy_496   :std_logic:='0';
  signal Energy_Bin_Rdy_497   :std_logic:='0';
  signal Energy_Bin_Rdy_498   :std_logic:='0';
  signal Energy_Bin_Rdy_499   :std_logic:='0';
  signal Energy_Bin_Rdy_500   :std_logic:='0';
  signal Energy_Bin_Rdy_501   :std_logic:='0';
  signal Energy_Bin_Rdy_502   :std_logic:='0';
  signal Energy_Bin_Rdy_503   :std_logic:='0';
  signal Energy_Bin_Rdy_504   :std_logic:='0';
  signal Energy_Bin_Rdy_505   :std_logic:='0';
  signal Energy_Bin_Rdy_506   :std_logic:='0';
  signal Energy_Bin_Rdy_507   :std_logic:='0';
  signal Energy_Bin_Rdy_508   :std_logic:='0';
  signal Energy_Bin_Rdy_509   :std_logic:='0';
  signal Energy_Bin_Rdy_510   :std_logic:='0';
  signal Energy_Bin_Rdy_511   :std_logic:='0';
  signal Energy_Bin_Rdy_512   :std_logic:='0';
  signal Energy_Bin_Rdy_513   :std_logic:='0';
  signal Energy_Bin_Rdy_514   :std_logic:='0';
  signal Energy_Bin_Rdy_515   :std_logic:='0';
  signal Energy_Bin_Rdy_516   :std_logic:='0';
  signal Energy_Bin_Rdy_517   :std_logic:='0';
  signal Energy_Bin_Rdy_518   :std_logic:='0';
  signal Energy_Bin_Rdy_519   :std_logic:='0';
  signal Energy_Bin_Rdy_520   :std_logic:='0';
  signal Energy_Bin_Rdy_521   :std_logic:='0';
  signal Energy_Bin_Rdy_522   :std_logic:='0';
  signal Energy_Bin_Rdy_523   :std_logic:='0';
  signal Energy_Bin_Rdy_524   :std_logic:='0';
  signal Energy_Bin_Rdy_525   :std_logic:='0';
  signal Energy_Bin_Rdy_526   :std_logic:='0';
  signal Energy_Bin_Rdy_527   :std_logic:='0';
  signal Energy_Bin_Rdy_528   :std_logic:='0';
  signal Energy_Bin_Rdy_529   :std_logic:='0';
  signal Energy_Bin_Rdy_530   :std_logic:='0';
  signal Energy_Bin_Rdy_531   :std_logic:='0';
  signal Energy_Bin_Rdy_532   :std_logic:='0';
  signal Energy_Bin_Rdy_533   :std_logic:='0';
  signal Energy_Bin_Rdy_534   :std_logic:='0';
  signal Energy_Bin_Rdy_535   :std_logic:='0';
  signal Energy_Bin_Rdy_536   :std_logic:='0';
  signal Energy_Bin_Rdy_537   :std_logic:='0';
  signal Energy_Bin_Rdy_538   :std_logic:='0';
  signal Energy_Bin_Rdy_539   :std_logic:='0';
  signal Energy_Bin_Rdy_540   :std_logic:='0';
  signal Energy_Bin_Rdy_541   :std_logic:='0';
  signal Energy_Bin_Rdy_542   :std_logic:='0';
  signal Energy_Bin_Rdy_543   :std_logic:='0';
  signal Energy_Bin_Rdy_544   :std_logic:='0';
  signal Energy_Bin_Rdy_545   :std_logic:='0';
  signal Energy_Bin_Rdy_546   :std_logic:='0';
  signal Energy_Bin_Rdy_547   :std_logic:='0';
  signal Energy_Bin_Rdy_548   :std_logic:='0';
  signal Energy_Bin_Rdy_549   :std_logic:='0';
  signal Energy_Bin_Rdy_550   :std_logic:='0';
  signal Energy_Bin_Rdy_551   :std_logic:='0';
  signal Energy_Bin_Rdy_552   :std_logic:='0';
  signal Energy_Bin_Rdy_553   :std_logic:='0';
  signal Energy_Bin_Rdy_554   :std_logic:='0';
  signal Energy_Bin_Rdy_555   :std_logic:='0';
  signal Energy_Bin_Rdy_556   :std_logic:='0';
  signal Energy_Bin_Rdy_557   :std_logic:='0';
  signal Energy_Bin_Rdy_558   :std_logic:='0';
  signal Energy_Bin_Rdy_559   :std_logic:='0';
  signal Energy_Bin_Rdy_560   :std_logic:='0';
  signal Energy_Bin_Rdy_561   :std_logic:='0';
  signal Energy_Bin_Rdy_562   :std_logic:='0';
  signal Energy_Bin_Rdy_563   :std_logic:='0';
  signal Energy_Bin_Rdy_564   :std_logic:='0';
  signal Energy_Bin_Rdy_565   :std_logic:='0';
  signal Energy_Bin_Rdy_566   :std_logic:='0';
  signal Energy_Bin_Rdy_567   :std_logic:='0';
  signal Energy_Bin_Rdy_568   :std_logic:='0';
  signal Energy_Bin_Rdy_569   :std_logic:='0';
  signal Energy_Bin_Rdy_570   :std_logic:='0';
  signal Energy_Bin_Rdy_571   :std_logic:='0';
  signal Energy_Bin_Rdy_572   :std_logic:='0';
  signal Energy_Bin_Rdy_573   :std_logic:='0';
  signal Energy_Bin_Rdy_574   :std_logic:='0';
  signal Energy_Bin_Rdy_575   :std_logic:='0';
  signal Energy_Bin_Rdy_576   :std_logic:='0';
  signal Energy_Bin_Rdy_577   :std_logic:='0';
  signal Energy_Bin_Rdy_578   :std_logic:='0';
  signal Energy_Bin_Rdy_579   :std_logic:='0';
  signal Energy_Bin_Rdy_580   :std_logic:='0';
  signal Energy_Bin_Rdy_581   :std_logic:='0';
  signal Energy_Bin_Rdy_582   :std_logic:='0';
  signal Energy_Bin_Rdy_583   :std_logic:='0';
  signal Energy_Bin_Rdy_584   :std_logic:='0';
  signal Energy_Bin_Rdy_585   :std_logic:='0';
  signal Energy_Bin_Rdy_586   :std_logic:='0';
  signal Energy_Bin_Rdy_587   :std_logic:='0';
  signal Energy_Bin_Rdy_588   :std_logic:='0';
  signal Energy_Bin_Rdy_589   :std_logic:='0';
  signal Energy_Bin_Rdy_590   :std_logic:='0';
  signal Energy_Bin_Rdy_591   :std_logic:='0';
  signal Energy_Bin_Rdy_592   :std_logic:='0';
  signal Energy_Bin_Rdy_593   :std_logic:='0';
  signal Energy_Bin_Rdy_594   :std_logic:='0';
  signal Energy_Bin_Rdy_595   :std_logic:='0';
  signal Energy_Bin_Rdy_596   :std_logic:='0';
  signal Energy_Bin_Rdy_597   :std_logic:='0';
  signal Energy_Bin_Rdy_598   :std_logic:='0';
  signal Energy_Bin_Rdy_599   :std_logic:='0';
  signal Energy_Bin_Rdy_600   :std_logic:='0';
  signal Energy_Bin_Rdy_601   :std_logic:='0';
  signal Energy_Bin_Rdy_602   :std_logic:='0';
  signal Energy_Bin_Rdy_603   :std_logic:='0';
  signal Energy_Bin_Rdy_604   :std_logic:='0';
  signal Energy_Bin_Rdy_605   :std_logic:='0';
  signal Energy_Bin_Rdy_606   :std_logic:='0';
  signal Energy_Bin_Rdy_607   :std_logic:='0';
  signal Energy_Bin_Rdy_608   :std_logic:='0';
  signal Energy_Bin_Rdy_609   :std_logic:='0';
  signal Energy_Bin_Rdy_610   :std_logic:='0';
  signal Energy_Bin_Rdy_611   :std_logic:='0';
  signal Energy_Bin_Rdy_612   :std_logic:='0';
  signal Energy_Bin_Rdy_613   :std_logic:='0';
  signal Energy_Bin_Rdy_614   :std_logic:='0';
  signal Energy_Bin_Rdy_615   :std_logic:='0';
  signal Energy_Bin_Rdy_616   :std_logic:='0';
  signal Energy_Bin_Rdy_617   :std_logic:='0';
  signal Energy_Bin_Rdy_618   :std_logic:='0';
  signal Energy_Bin_Rdy_619   :std_logic:='0';
  signal Energy_Bin_Rdy_620   :std_logic:='0';
  signal Energy_Bin_Rdy_621   :std_logic:='0';
  signal Energy_Bin_Rdy_622   :std_logic:='0';
  signal Energy_Bin_Rdy_623   :std_logic:='0';
  signal Energy_Bin_Rdy_624   :std_logic:='0';
  signal Energy_Bin_Rdy_625   :std_logic:='0';
  signal Energy_Bin_Rdy_626   :std_logic:='0';
  signal Energy_Bin_Rdy_627   :std_logic:='0';
  signal Energy_Bin_Rdy_628   :std_logic:='0';
  signal Energy_Bin_Rdy_629   :std_logic:='0';
  signal Energy_Bin_Rdy_630   :std_logic:='0';
  signal Energy_Bin_Rdy_631   :std_logic:='0';
  signal Energy_Bin_Rdy_632   :std_logic:='0';
  signal Energy_Bin_Rdy_633   :std_logic:='0';
  signal Energy_Bin_Rdy_634   :std_logic:='0';
  signal Energy_Bin_Rdy_635   :std_logic:='0';
  signal Energy_Bin_Rdy_636   :std_logic:='0';
  signal Energy_Bin_Rdy_637   :std_logic:='0';
  signal Energy_Bin_Rdy_638   :std_logic:='0';
  signal Energy_Bin_Rdy_639   :std_logic:='0';
  signal Energy_Bin_Rdy_640   :std_logic:='0';
  signal Energy_Bin_Rdy_641   :std_logic:='0';
  signal Energy_Bin_Rdy_642   :std_logic:='0';
  signal Energy_Bin_Rdy_643   :std_logic:='0';
  signal Energy_Bin_Rdy_644   :std_logic:='0';
  signal Energy_Bin_Rdy_645   :std_logic:='0';
  signal Energy_Bin_Rdy_646   :std_logic:='0';
  signal Energy_Bin_Rdy_647   :std_logic:='0';
  signal Energy_Bin_Rdy_648   :std_logic:='0';
  signal Energy_Bin_Rdy_649   :std_logic:='0';
  signal Energy_Bin_Rdy_650   :std_logic:='0';
  signal Energy_Bin_Rdy_651   :std_logic:='0';
  signal Energy_Bin_Rdy_652   :std_logic:='0';
  signal Energy_Bin_Rdy_653   :std_logic:='0';
  signal Energy_Bin_Rdy_654   :std_logic:='0';
  signal Energy_Bin_Rdy_655   :std_logic:='0';
  signal Energy_Bin_Rdy_656   :std_logic:='0';
  signal Energy_Bin_Rdy_657   :std_logic:='0';
  signal Energy_Bin_Rdy_658   :std_logic:='0';
  signal Energy_Bin_Rdy_659   :std_logic:='0';
  signal Energy_Bin_Rdy_660   :std_logic:='0';
  signal Energy_Bin_Rdy_661   :std_logic:='0';
  signal Energy_Bin_Rdy_662   :std_logic:='0';
  signal Energy_Bin_Rdy_663   :std_logic:='0';
  signal Energy_Bin_Rdy_664   :std_logic:='0';
  signal Energy_Bin_Rdy_665   :std_logic:='0';
  signal Energy_Bin_Rdy_666   :std_logic:='0';
  signal Energy_Bin_Rdy_667   :std_logic:='0';
  signal Energy_Bin_Rdy_668   :std_logic:='0';
  signal Energy_Bin_Rdy_669   :std_logic:='0';
  signal Energy_Bin_Rdy_670   :std_logic:='0';
  signal Energy_Bin_Rdy_671   :std_logic:='0';
  signal Energy_Bin_Rdy_672   :std_logic:='0';
  signal Energy_Bin_Rdy_673   :std_logic:='0';
  signal Energy_Bin_Rdy_674   :std_logic:='0';
  signal Energy_Bin_Rdy_675   :std_logic:='0';
  signal Energy_Bin_Rdy_676   :std_logic:='0';
  signal Energy_Bin_Rdy_677   :std_logic:='0';
  signal Energy_Bin_Rdy_678   :std_logic:='0';
  signal Energy_Bin_Rdy_679   :std_logic:='0';
  signal Energy_Bin_Rdy_680   :std_logic:='0';
  signal Energy_Bin_Rdy_681   :std_logic:='0';
  signal Energy_Bin_Rdy_682   :std_logic:='0';
  signal Energy_Bin_Rdy_683   :std_logic:='0';
  signal Energy_Bin_Rdy_684   :std_logic:='0';
  signal Energy_Bin_Rdy_685   :std_logic:='0';
  signal Energy_Bin_Rdy_686   :std_logic:='0';
  signal Energy_Bin_Rdy_687   :std_logic:='0';
  signal Energy_Bin_Rdy_688   :std_logic:='0';
  signal Energy_Bin_Rdy_689   :std_logic:='0';
  signal Energy_Bin_Rdy_690   :std_logic:='0';
  signal Energy_Bin_Rdy_691   :std_logic:='0';
  signal Energy_Bin_Rdy_692   :std_logic:='0';
  signal Energy_Bin_Rdy_693   :std_logic:='0';
  signal Energy_Bin_Rdy_694   :std_logic:='0';
  signal Energy_Bin_Rdy_695   :std_logic:='0';
  signal Energy_Bin_Rdy_696   :std_logic:='0';
  signal Energy_Bin_Rdy_697   :std_logic:='0';
  signal Energy_Bin_Rdy_698   :std_logic:='0';
  signal Energy_Bin_Rdy_699   :std_logic:='0';
  signal Energy_Bin_Rdy_700   :std_logic:='0';
  signal Energy_Bin_Rdy_701   :std_logic:='0';
  signal Energy_Bin_Rdy_702   :std_logic:='0';
  signal Energy_Bin_Rdy_703   :std_logic:='0';
  signal Energy_Bin_Rdy_704   :std_logic:='0';
  signal Energy_Bin_Rdy_705   :std_logic:='0';
  signal Energy_Bin_Rdy_706   :std_logic:='0';
  signal Energy_Bin_Rdy_707   :std_logic:='0';
  signal Energy_Bin_Rdy_708   :std_logic:='0';
  signal Energy_Bin_Rdy_709   :std_logic:='0';
  signal Energy_Bin_Rdy_710   :std_logic:='0';
  signal Energy_Bin_Rdy_711   :std_logic:='0';
  signal Energy_Bin_Rdy_712   :std_logic:='0';
  signal Energy_Bin_Rdy_713   :std_logic:='0';
  signal Energy_Bin_Rdy_714   :std_logic:='0';
  signal Energy_Bin_Rdy_715   :std_logic:='0';
  signal Energy_Bin_Rdy_716   :std_logic:='0';
  signal Energy_Bin_Rdy_717   :std_logic:='0';
  signal Energy_Bin_Rdy_718   :std_logic:='0';
  signal Energy_Bin_Rdy_719   :std_logic:='0';
  signal Energy_Bin_Rdy_720   :std_logic:='0';
  signal Energy_Bin_Rdy_721   :std_logic:='0';
  signal Energy_Bin_Rdy_722   :std_logic:='0';
  signal Energy_Bin_Rdy_723   :std_logic:='0';
  signal Energy_Bin_Rdy_724   :std_logic:='0';
  signal Energy_Bin_Rdy_725   :std_logic:='0';
  signal Energy_Bin_Rdy_726   :std_logic:='0';
  signal Energy_Bin_Rdy_727   :std_logic:='0';
  signal Energy_Bin_Rdy_728   :std_logic:='0';
  signal Energy_Bin_Rdy_729   :std_logic:='0';
  signal Energy_Bin_Rdy_730   :std_logic:='0';
  signal Energy_Bin_Rdy_731   :std_logic:='0';
  signal Energy_Bin_Rdy_732   :std_logic:='0';
  signal Energy_Bin_Rdy_733   :std_logic:='0';
  signal Energy_Bin_Rdy_734   :std_logic:='0';
  signal Energy_Bin_Rdy_735   :std_logic:='0';
  signal Energy_Bin_Rdy_736   :std_logic:='0';
  signal Energy_Bin_Rdy_737   :std_logic:='0';
  signal Energy_Bin_Rdy_738   :std_logic:='0';
  signal Energy_Bin_Rdy_739   :std_logic:='0';
  signal Energy_Bin_Rdy_740   :std_logic:='0';
  signal Energy_Bin_Rdy_741   :std_logic:='0';
  signal Energy_Bin_Rdy_742   :std_logic:='0';
  signal Energy_Bin_Rdy_743   :std_logic:='0';
  signal Energy_Bin_Rdy_744   :std_logic:='0';
  signal Energy_Bin_Rdy_745   :std_logic:='0';
  signal Energy_Bin_Rdy_746   :std_logic:='0';
  signal Energy_Bin_Rdy_747   :std_logic:='0';
  signal Energy_Bin_Rdy_748   :std_logic:='0';
  signal Energy_Bin_Rdy_749   :std_logic:='0';
  signal Energy_Bin_Rdy_750   :std_logic:='0';
  signal Energy_Bin_Rdy_751   :std_logic:='0';
  signal Energy_Bin_Rdy_752   :std_logic:='0';
  signal Energy_Bin_Rdy_753   :std_logic:='0';
  signal Energy_Bin_Rdy_754   :std_logic:='0';
  signal Energy_Bin_Rdy_755   :std_logic:='0';
  signal Energy_Bin_Rdy_756   :std_logic:='0';
  signal Energy_Bin_Rdy_757   :std_logic:='0';
  signal Energy_Bin_Rdy_758   :std_logic:='0';
  signal Energy_Bin_Rdy_759   :std_logic:='0';
  signal Energy_Bin_Rdy_760   :std_logic:='0';
  signal Energy_Bin_Rdy_761   :std_logic:='0';
  signal Energy_Bin_Rdy_762   :std_logic:='0';
  signal Energy_Bin_Rdy_763   :std_logic:='0';
  signal Energy_Bin_Rdy_764   :std_logic:='0';
  signal Energy_Bin_Rdy_765   :std_logic:='0';
  signal Energy_Bin_Rdy_766   :std_logic:='0';
  signal Energy_Bin_Rdy_767   :std_logic:='0';
  signal Energy_Bin_Rdy_768   :std_logic:='0';
  signal Energy_Bin_Rdy_769   :std_logic:='0';
  signal Energy_Bin_Rdy_770   :std_logic:='0';
  signal Energy_Bin_Rdy_771   :std_logic:='0';
  signal Energy_Bin_Rdy_772   :std_logic:='0';
  signal Energy_Bin_Rdy_773   :std_logic:='0';
  signal Energy_Bin_Rdy_774   :std_logic:='0';
  signal Energy_Bin_Rdy_775   :std_logic:='0';
  signal Energy_Bin_Rdy_776   :std_logic:='0';
  signal Energy_Bin_Rdy_777   :std_logic:='0';
  signal Energy_Bin_Rdy_778   :std_logic:='0';
  signal Energy_Bin_Rdy_779   :std_logic:='0';
  signal Energy_Bin_Rdy_780   :std_logic:='0';
  signal Energy_Bin_Rdy_781   :std_logic:='0';
  signal Energy_Bin_Rdy_782   :std_logic:='0';
  signal Energy_Bin_Rdy_783   :std_logic:='0';
  signal Energy_Bin_Rdy_784   :std_logic:='0';
  signal Energy_Bin_Rdy_785   :std_logic:='0';
  signal Energy_Bin_Rdy_786   :std_logic:='0';
  signal Energy_Bin_Rdy_787   :std_logic:='0';
  signal Energy_Bin_Rdy_788   :std_logic:='0';
  signal Energy_Bin_Rdy_789   :std_logic:='0';
  signal Energy_Bin_Rdy_790   :std_logic:='0';
  signal Energy_Bin_Rdy_791   :std_logic:='0';
  signal Energy_Bin_Rdy_792   :std_logic:='0';
  signal Energy_Bin_Rdy_793   :std_logic:='0';
  signal Energy_Bin_Rdy_794   :std_logic:='0';
  signal Energy_Bin_Rdy_795   :std_logic:='0';
  signal Energy_Bin_Rdy_796   :std_logic:='0';
  signal Energy_Bin_Rdy_797   :std_logic:='0';
  signal Energy_Bin_Rdy_798   :std_logic:='0';
  signal Energy_Bin_Rdy_799   :std_logic:='0';
  signal Energy_Bin_Rdy_800   :std_logic:='0';
  signal Energy_Bin_Rdy_801   :std_logic:='0';
  signal Energy_Bin_Rdy_802   :std_logic:='0';
  signal Energy_Bin_Rdy_803   :std_logic:='0';
  signal Energy_Bin_Rdy_804   :std_logic:='0';
  signal Energy_Bin_Rdy_805   :std_logic:='0';
  signal Energy_Bin_Rdy_806   :std_logic:='0';
  signal Energy_Bin_Rdy_807   :std_logic:='0';
  signal Energy_Bin_Rdy_808   :std_logic:='0';
  signal Energy_Bin_Rdy_809   :std_logic:='0';
  signal Energy_Bin_Rdy_810   :std_logic:='0';
  signal Energy_Bin_Rdy_811   :std_logic:='0';
  signal Energy_Bin_Rdy_812   :std_logic:='0';
  signal Energy_Bin_Rdy_813   :std_logic:='0';
  signal Energy_Bin_Rdy_814   :std_logic:='0';
  signal Energy_Bin_Rdy_815   :std_logic:='0';
  signal Energy_Bin_Rdy_816   :std_logic:='0';
  signal Energy_Bin_Rdy_817   :std_logic:='0';
  signal Energy_Bin_Rdy_818   :std_logic:='0';
  signal Energy_Bin_Rdy_819   :std_logic:='0';
  signal Energy_Bin_Rdy_820   :std_logic:='0';
  signal Energy_Bin_Rdy_821   :std_logic:='0';
  signal Energy_Bin_Rdy_822   :std_logic:='0';
  signal Energy_Bin_Rdy_823   :std_logic:='0';
  signal Energy_Bin_Rdy_824   :std_logic:='0';
  signal Energy_Bin_Rdy_825   :std_logic:='0';
  signal Energy_Bin_Rdy_826   :std_logic:='0';
  signal Energy_Bin_Rdy_827   :std_logic:='0';
  signal Energy_Bin_Rdy_828   :std_logic:='0';
  signal Energy_Bin_Rdy_829   :std_logic:='0';
  signal Energy_Bin_Rdy_830   :std_logic:='0';
  signal Energy_Bin_Rdy_831   :std_logic:='0';
  signal Energy_Bin_Rdy_832   :std_logic:='0';
  signal Energy_Bin_Rdy_833   :std_logic:='0';
  signal Energy_Bin_Rdy_834   :std_logic:='0';
  signal Energy_Bin_Rdy_835   :std_logic:='0';
  signal Energy_Bin_Rdy_836   :std_logic:='0';
  signal Energy_Bin_Rdy_837   :std_logic:='0';
  signal Energy_Bin_Rdy_838   :std_logic:='0';
  signal Energy_Bin_Rdy_839   :std_logic:='0';
  signal Energy_Bin_Rdy_840   :std_logic:='0';
  signal Energy_Bin_Rdy_841   :std_logic:='0';
  signal Energy_Bin_Rdy_842   :std_logic:='0';
  signal Energy_Bin_Rdy_843   :std_logic:='0';
  signal Energy_Bin_Rdy_844   :std_logic:='0';
  signal Energy_Bin_Rdy_845   :std_logic:='0';
  signal Energy_Bin_Rdy_846   :std_logic:='0';
  signal Energy_Bin_Rdy_847   :std_logic:='0';
  signal Energy_Bin_Rdy_848   :std_logic:='0';
  signal Energy_Bin_Rdy_849   :std_logic:='0';
  signal Energy_Bin_Rdy_850   :std_logic:='0';
  signal Energy_Bin_Rdy_851   :std_logic:='0';
  signal Energy_Bin_Rdy_852   :std_logic:='0';
  signal Energy_Bin_Rdy_853   :std_logic:='0';
  signal Energy_Bin_Rdy_854   :std_logic:='0';
  signal Energy_Bin_Rdy_855   :std_logic:='0';
  signal Energy_Bin_Rdy_856   :std_logic:='0';
  signal Energy_Bin_Rdy_857   :std_logic:='0';
  signal Energy_Bin_Rdy_858   :std_logic:='0';
  signal Energy_Bin_Rdy_859   :std_logic:='0';
  signal Energy_Bin_Rdy_860   :std_logic:='0';
  signal Energy_Bin_Rdy_861   :std_logic:='0';
  signal Energy_Bin_Rdy_862   :std_logic:='0';
  signal Energy_Bin_Rdy_863   :std_logic:='0';
  signal Energy_Bin_Rdy_864   :std_logic:='0';
  signal Energy_Bin_Rdy_865   :std_logic:='0';
  signal Energy_Bin_Rdy_866   :std_logic:='0';
  signal Energy_Bin_Rdy_867   :std_logic:='0';
  signal Energy_Bin_Rdy_868   :std_logic:='0';
  signal Energy_Bin_Rdy_869   :std_logic:='0';
  signal Energy_Bin_Rdy_870   :std_logic:='0';
  signal Energy_Bin_Rdy_871   :std_logic:='0';
  signal Energy_Bin_Rdy_872   :std_logic:='0';
  signal Energy_Bin_Rdy_873   :std_logic:='0';
  signal Energy_Bin_Rdy_874   :std_logic:='0';
  signal Energy_Bin_Rdy_875   :std_logic:='0';
  signal Energy_Bin_Rdy_876   :std_logic:='0';
  signal Energy_Bin_Rdy_877   :std_logic:='0';
  signal Energy_Bin_Rdy_878   :std_logic:='0';
  signal Energy_Bin_Rdy_879   :std_logic:='0';
  signal Energy_Bin_Rdy_880   :std_logic:='0';
  signal Energy_Bin_Rdy_881   :std_logic:='0';
  signal Energy_Bin_Rdy_882   :std_logic:='0';
  signal Energy_Bin_Rdy_883   :std_logic:='0';
  signal Energy_Bin_Rdy_884   :std_logic:='0';
  signal Energy_Bin_Rdy_885   :std_logic:='0';
  signal Energy_Bin_Rdy_886   :std_logic:='0';
  signal Energy_Bin_Rdy_887   :std_logic:='0';
  signal Energy_Bin_Rdy_888   :std_logic:='0';
  signal Energy_Bin_Rdy_889   :std_logic:='0';
  signal Energy_Bin_Rdy_890   :std_logic:='0';
  signal Energy_Bin_Rdy_891   :std_logic:='0';
  signal Energy_Bin_Rdy_892   :std_logic:='0';
  signal Energy_Bin_Rdy_893   :std_logic:='0';
  signal Energy_Bin_Rdy_894   :std_logic:='0';
  signal Energy_Bin_Rdy_895   :std_logic:='0';
  signal Energy_Bin_Rdy_896   :std_logic:='0';
  signal Energy_Bin_Rdy_897   :std_logic:='0';
  signal Energy_Bin_Rdy_898   :std_logic:='0';
  signal Energy_Bin_Rdy_899   :std_logic:='0';
  signal Energy_Bin_Rdy_900   :std_logic:='0';
  signal Energy_Bin_Rdy_901   :std_logic:='0';
  signal Energy_Bin_Rdy_902   :std_logic:='0';
  signal Energy_Bin_Rdy_903   :std_logic:='0';
  signal Energy_Bin_Rdy_904   :std_logic:='0';
  signal Energy_Bin_Rdy_905   :std_logic:='0';
  signal Energy_Bin_Rdy_906   :std_logic:='0';
  signal Energy_Bin_Rdy_907   :std_logic:='0';
  signal Energy_Bin_Rdy_908   :std_logic:='0';
  signal Energy_Bin_Rdy_909   :std_logic:='0';
  signal Energy_Bin_Rdy_910   :std_logic:='0';
  signal Energy_Bin_Rdy_911   :std_logic:='0';
  signal Energy_Bin_Rdy_912   :std_logic:='0';
  signal Energy_Bin_Rdy_913   :std_logic:='0';
  signal Energy_Bin_Rdy_914   :std_logic:='0';
  signal Energy_Bin_Rdy_915   :std_logic:='0';
  signal Energy_Bin_Rdy_916   :std_logic:='0';
  signal Energy_Bin_Rdy_917   :std_logic:='0';
  signal Energy_Bin_Rdy_918   :std_logic:='0';
  signal Energy_Bin_Rdy_919   :std_logic:='0';
  signal Energy_Bin_Rdy_920   :std_logic:='0';
  signal Energy_Bin_Rdy_921   :std_logic:='0';
  signal Energy_Bin_Rdy_922   :std_logic:='0';
  signal Energy_Bin_Rdy_923   :std_logic:='0';
  signal Energy_Bin_Rdy_924   :std_logic:='0';
  signal Energy_Bin_Rdy_925   :std_logic:='0';
  signal Energy_Bin_Rdy_926   :std_logic:='0';
  signal Energy_Bin_Rdy_927   :std_logic:='0';
  signal Energy_Bin_Rdy_928   :std_logic:='0';
  signal Energy_Bin_Rdy_929   :std_logic:='0';
  signal Energy_Bin_Rdy_930   :std_logic:='0';
  signal Energy_Bin_Rdy_931   :std_logic:='0';
  signal Energy_Bin_Rdy_932   :std_logic:='0';
  signal Energy_Bin_Rdy_933   :std_logic:='0';
  signal Energy_Bin_Rdy_934   :std_logic:='0';
  signal Energy_Bin_Rdy_935   :std_logic:='0';
  signal Energy_Bin_Rdy_936   :std_logic:='0';
  signal Energy_Bin_Rdy_937   :std_logic:='0';
  signal Energy_Bin_Rdy_938   :std_logic:='0';
  signal Energy_Bin_Rdy_939   :std_logic:='0';
  signal Energy_Bin_Rdy_940   :std_logic:='0';
  signal Energy_Bin_Rdy_941   :std_logic:='0';
  signal Energy_Bin_Rdy_942   :std_logic:='0';
  signal Energy_Bin_Rdy_943   :std_logic:='0';
  signal Energy_Bin_Rdy_944   :std_logic:='0';
  signal Energy_Bin_Rdy_945   :std_logic:='0';
  signal Energy_Bin_Rdy_946   :std_logic:='0';
  signal Energy_Bin_Rdy_947   :std_logic:='0';
  signal Energy_Bin_Rdy_948   :std_logic:='0';
  signal Energy_Bin_Rdy_949   :std_logic:='0';
  signal Energy_Bin_Rdy_950   :std_logic:='0';
  signal Energy_Bin_Rdy_951   :std_logic:='0';
  signal Energy_Bin_Rdy_952   :std_logic:='0';
  signal Energy_Bin_Rdy_953   :std_logic:='0';
  signal Energy_Bin_Rdy_954   :std_logic:='0';
  signal Energy_Bin_Rdy_955   :std_logic:='0';
  signal Energy_Bin_Rdy_956   :std_logic:='0';
  signal Energy_Bin_Rdy_957   :std_logic:='0';
  signal Energy_Bin_Rdy_958   :std_logic:='0';
  signal Energy_Bin_Rdy_959   :std_logic:='0';
  signal Energy_Bin_Rdy_960   :std_logic:='0';
  signal Energy_Bin_Rdy_961   :std_logic:='0';
  signal Energy_Bin_Rdy_962   :std_logic:='0';
  signal Energy_Bin_Rdy_963   :std_logic:='0';
  signal Energy_Bin_Rdy_964   :std_logic:='0';
  signal Energy_Bin_Rdy_965   :std_logic:='0';
  signal Energy_Bin_Rdy_966   :std_logic:='0';
  signal Energy_Bin_Rdy_967   :std_logic:='0';
  signal Energy_Bin_Rdy_968   :std_logic:='0';
  signal Energy_Bin_Rdy_969   :std_logic:='0';
  signal Energy_Bin_Rdy_970   :std_logic:='0';
  signal Energy_Bin_Rdy_971   :std_logic:='0';
  signal Energy_Bin_Rdy_972   :std_logic:='0';
  signal Energy_Bin_Rdy_973   :std_logic:='0';
  signal Energy_Bin_Rdy_974   :std_logic:='0';
  signal Energy_Bin_Rdy_975   :std_logic:='0';
  signal Energy_Bin_Rdy_976   :std_logic:='0';
  signal Energy_Bin_Rdy_977   :std_logic:='0';
  signal Energy_Bin_Rdy_978   :std_logic:='0';
  signal Energy_Bin_Rdy_979   :std_logic:='0';
  signal Energy_Bin_Rdy_980   :std_logic:='0';
  signal Energy_Bin_Rdy_981   :std_logic:='0';
  signal Energy_Bin_Rdy_982   :std_logic:='0';
  signal Energy_Bin_Rdy_983   :std_logic:='0';
  signal Energy_Bin_Rdy_984   :std_logic:='0';
  signal Energy_Bin_Rdy_985   :std_logic:='0';
  signal Energy_Bin_Rdy_986   :std_logic:='0';
  signal Energy_Bin_Rdy_987   :std_logic:='0';
  signal Energy_Bin_Rdy_988   :std_logic:='0';
  signal Energy_Bin_Rdy_989   :std_logic:='0';
  signal Energy_Bin_Rdy_990   :std_logic:='0';
  signal Energy_Bin_Rdy_991   :std_logic:='0';
  signal Energy_Bin_Rdy_992   :std_logic:='0';
  signal Energy_Bin_Rdy_993   :std_logic:='0';
  signal Energy_Bin_Rdy_994   :std_logic:='0';
  signal Energy_Bin_Rdy_995   :std_logic:='0';
  signal Energy_Bin_Rdy_996   :std_logic:='0';
  signal Energy_Bin_Rdy_997   :std_logic:='0';
  signal Energy_Bin_Rdy_998   :std_logic:='0';
  signal Energy_Bin_Rdy_999   :std_logic:='0';
  signal Energy_Bin_Rdy_1000  :std_logic:='0';
  signal Energy_Bin_Rdy_1001  :std_logic:='0';
  signal Energy_Bin_Rdy_1002  :std_logic:='0';
  signal Energy_Bin_Rdy_1003  :std_logic:='0';
  signal Energy_Bin_Rdy_1004  :std_logic:='0';
  signal Energy_Bin_Rdy_1005  :std_logic:='0';
  signal Energy_Bin_Rdy_1006  :std_logic:='0';
  signal Energy_Bin_Rdy_1007  :std_logic:='0';
  signal Energy_Bin_Rdy_1008  :std_logic:='0';
  signal Energy_Bin_Rdy_1009  :std_logic:='0';
  signal Energy_Bin_Rdy_1010  :std_logic:='0';
  signal Energy_Bin_Rdy_1011  :std_logic:='0';
  signal Energy_Bin_Rdy_1012  :std_logic:='0';
  signal Energy_Bin_Rdy_1013  :std_logic:='0';
  signal Energy_Bin_Rdy_1014  :std_logic:='0';
  signal Energy_Bin_Rdy_1015  :std_logic:='0';
  signal Energy_Bin_Rdy_1016  :std_logic:='0';
  signal Energy_Bin_Rdy_1017  :std_logic:='0';
  signal Energy_Bin_Rdy_1018  :std_logic:='0';
  signal Energy_Bin_Rdy_1019  :std_logic:='0';
  signal Energy_Bin_Rdy_1020  :std_logic:='0';
  signal Energy_Bin_Rdy_1021  :std_logic:='0';
  signal Energy_Bin_Rdy_1022  :std_logic:='0';
  signal Energy_Bin_Rdy_1023  :std_logic:='0';
  signal Energy_Bin_Rdy_1024  :std_logic:='0';
  
  signal PEAK_FL_C1       			 :std_logic:='0'; /* synthesis preserve=1*/
  signal PEAK_FL_C1_s1    			 :std_logic:='0'; /* synthesis preserve=1*/
  signal PEAK_FL_C1_s2    			 :std_logic:='0'; /* synthesis preserve=1*/
  signal PEAK_FL_Ris      			 :std_logic:='0'; /* synthesis preserve=1*/
  signal PEAK_FL_Ris_s    			 :std_logic:='0'; /* synthesis preserve=1*/
  signal Energy_Ris_Dis   			 :std_logic:='0'; /* synthesis preserve=1*/

  signal PEAK_FL_C1_pos       		 :std_logic:='0'; /* synthesis preserve=1*/
  signal PEAK_FL_C1_pos_s1    		 :std_logic:='0'; /* synthesis preserve=1*/
  signal PEAK_FL_C1_pos_s2    		 :std_logic:='0'; /* synthesis preserve=1*/
  signal PEAK_FL_Ris_pos      		 :std_logic:='0'; /* synthesis preserve=1*/
  signal PEAK_FL_Ris_pos_s    		 :std_logic:='0'; /* synthesis preserve=1*/
  signal Energy_Ris_Dis_pos   		 :std_logic:='0'; /* synthesis preserve=1*/
  
  signal s_Energy_Bin_reject         :std_logic_vector(15 downto 0); 
  signal s_Energy_Bin_Pos_reject     :std_logic_vector(15 downto 0);
  signal Energy_Bin_Pos_rdy          :std_logic;
  signal Energy_Bin_Pos_rdy_reject   :std_logic;
  signal Energy_Bin_rdy_reject       :std_logic;


  signal Bin_OR		          		 :std_logic:='0';  
  signal Bin_OR_pos          		 :std_logic:='0'; 
  
  signal wr_cnt           :std_logic_vector(31 downto 0)
                          :=(others =>'0');  		                                          
                     	                                                   
--+----------
-- Start of architecture code
--+----------
begin
  --+----------
  -- Global signal assignments for the architecture.
  --+----------

  o_Energy_Bin_Pos_1    <= s_Energy_Bin_Pos_1    ;
  o_Energy_Bin_Pos_2    <= s_Energy_Bin_Pos_2    ;
  o_Energy_Bin_Pos_3    <= s_Energy_Bin_Pos_3    ;
  o_Energy_Bin_Pos_4    <= s_Energy_Bin_Pos_4    ;
  o_Energy_Bin_Pos_5    <= s_Energy_Bin_Pos_5    ;
  o_Energy_Bin_Pos_6    <= s_Energy_Bin_Pos_6    ;
  o_Energy_Bin_Pos_7    <= s_Energy_Bin_Pos_7    ;
  o_Energy_Bin_Pos_8    <= s_Energy_Bin_Pos_8    ;
  o_Energy_Bin_Pos_9    <= s_Energy_Bin_Pos_9    ;
  o_Energy_Bin_Pos_10   <= s_Energy_Bin_Pos_10   ;
  o_Energy_Bin_Pos_11   <= s_Energy_Bin_Pos_11   ;
  o_Energy_Bin_Pos_12   <= s_Energy_Bin_Pos_12   ;
  o_Energy_Bin_Pos_13   <= s_Energy_Bin_Pos_13   ;
  o_Energy_Bin_Pos_14   <= s_Energy_Bin_Pos_14   ;
  o_Energy_Bin_Pos_15   <= s_Energy_Bin_Pos_15   ;
  o_Energy_Bin_Pos_16   <= s_Energy_Bin_Pos_16   ;
  o_Energy_Bin_Pos_17   <= s_Energy_Bin_Pos_17   ;
  o_Energy_Bin_Pos_18   <= s_Energy_Bin_Pos_18   ;
  o_Energy_Bin_Pos_19   <= s_Energy_Bin_Pos_19   ;
  o_Energy_Bin_Pos_20   <= s_Energy_Bin_Pos_20   ;
  o_Energy_Bin_Pos_21   <= s_Energy_Bin_Pos_21   ;
  o_Energy_Bin_Pos_22   <= s_Energy_Bin_Pos_22   ;
  o_Energy_Bin_Pos_23   <= s_Energy_Bin_Pos_23   ;
  o_Energy_Bin_Pos_24   <= s_Energy_Bin_Pos_24   ;
  o_Energy_Bin_Pos_25   <= s_Energy_Bin_Pos_25   ;
  o_Energy_Bin_Pos_26   <= s_Energy_Bin_Pos_26   ;
  o_Energy_Bin_Pos_27   <= s_Energy_Bin_Pos_27   ;
  o_Energy_Bin_Pos_28   <= s_Energy_Bin_Pos_28   ;
  o_Energy_Bin_Pos_29   <= s_Energy_Bin_Pos_29   ;
  o_Energy_Bin_Pos_30   <= s_Energy_Bin_Pos_30   ;
  o_Energy_Bin_Pos_31   <= s_Energy_Bin_Pos_31   ;
  o_Energy_Bin_Pos_32   <= s_Energy_Bin_Pos_32   ;
  o_Energy_Bin_Pos_33   <= s_Energy_Bin_Pos_33   ;
  o_Energy_Bin_Pos_34   <= s_Energy_Bin_Pos_34   ;
  o_Energy_Bin_Pos_35   <= s_Energy_Bin_Pos_35   ;
  o_Energy_Bin_Pos_36   <= s_Energy_Bin_Pos_36   ;
  o_Energy_Bin_Pos_37   <= s_Energy_Bin_Pos_37   ;
  o_Energy_Bin_Pos_38   <= s_Energy_Bin_Pos_38   ;
  o_Energy_Bin_Pos_39   <= s_Energy_Bin_Pos_39   ;
  o_Energy_Bin_Pos_40   <= s_Energy_Bin_Pos_40   ;
  o_Energy_Bin_Pos_41   <= s_Energy_Bin_Pos_41   ;
  o_Energy_Bin_Pos_42   <= s_Energy_Bin_Pos_42   ;
  o_Energy_Bin_Pos_43   <= s_Energy_Bin_Pos_43   ;
  o_Energy_Bin_Pos_44   <= s_Energy_Bin_Pos_44   ;
  o_Energy_Bin_Pos_45   <= s_Energy_Bin_Pos_45   ;
  o_Energy_Bin_Pos_46   <= s_Energy_Bin_Pos_46   ;
  o_Energy_Bin_Pos_47   <= s_Energy_Bin_Pos_47   ;
  o_Energy_Bin_Pos_48   <= s_Energy_Bin_Pos_48   ;
  o_Energy_Bin_Pos_49   <= s_Energy_Bin_Pos_49   ;
  o_Energy_Bin_Pos_50   <= s_Energy_Bin_Pos_50   ;
  o_Energy_Bin_Pos_51   <= s_Energy_Bin_Pos_51   ;
  o_Energy_Bin_Pos_52   <= s_Energy_Bin_Pos_52   ;
  o_Energy_Bin_Pos_53   <= s_Energy_Bin_Pos_53   ;
  o_Energy_Bin_Pos_54   <= s_Energy_Bin_Pos_54   ;
  o_Energy_Bin_Pos_55   <= s_Energy_Bin_Pos_55   ;
  o_Energy_Bin_Pos_56   <= s_Energy_Bin_Pos_56   ;
  o_Energy_Bin_Pos_57   <= s_Energy_Bin_Pos_57   ;
  o_Energy_Bin_Pos_58   <= s_Energy_Bin_Pos_58   ;
  o_Energy_Bin_Pos_59   <= s_Energy_Bin_Pos_59   ;
  o_Energy_Bin_Pos_60   <= s_Energy_Bin_Pos_60   ;
  o_Energy_Bin_Pos_61   <= s_Energy_Bin_Pos_61   ;
  o_Energy_Bin_Pos_62   <= s_Energy_Bin_Pos_62   ;
  o_Energy_Bin_Pos_63   <= s_Energy_Bin_Pos_63   ;
  o_Energy_Bin_Pos_64   <= s_Energy_Bin_Pos_64   ;
  o_Energy_Bin_Pos_65   <= s_Energy_Bin_Pos_65   ;
  o_Energy_Bin_Pos_66   <= s_Energy_Bin_Pos_66   ;
  o_Energy_Bin_Pos_67   <= s_Energy_Bin_Pos_67   ;
  o_Energy_Bin_Pos_68   <= s_Energy_Bin_Pos_68   ;
  o_Energy_Bin_Pos_69   <= s_Energy_Bin_Pos_69   ;
  o_Energy_Bin_Pos_70   <= s_Energy_Bin_Pos_70   ;
  o_Energy_Bin_Pos_71   <= s_Energy_Bin_Pos_71   ;
  o_Energy_Bin_Pos_72   <= s_Energy_Bin_Pos_72   ;
  o_Energy_Bin_Pos_73   <= s_Energy_Bin_Pos_73   ;
  o_Energy_Bin_Pos_74   <= s_Energy_Bin_Pos_74   ;
  o_Energy_Bin_Pos_75   <= s_Energy_Bin_Pos_75   ;
  o_Energy_Bin_Pos_76   <= s_Energy_Bin_Pos_76   ;
  o_Energy_Bin_Pos_77   <= s_Energy_Bin_Pos_77   ;
  o_Energy_Bin_Pos_78   <= s_Energy_Bin_Pos_78   ;
  o_Energy_Bin_Pos_79   <= s_Energy_Bin_Pos_79   ;
  o_Energy_Bin_Pos_80   <= s_Energy_Bin_Pos_80   ;
  o_Energy_Bin_Pos_81   <= s_Energy_Bin_Pos_81   ;
  o_Energy_Bin_Pos_82   <= s_Energy_Bin_Pos_82   ;
  o_Energy_Bin_Pos_83   <= s_Energy_Bin_Pos_83   ;
  o_Energy_Bin_Pos_84   <= s_Energy_Bin_Pos_84   ;
  o_Energy_Bin_Pos_85   <= s_Energy_Bin_Pos_85   ;
  o_Energy_Bin_Pos_86   <= s_Energy_Bin_Pos_86   ;
  o_Energy_Bin_Pos_87   <= s_Energy_Bin_Pos_87   ;
  o_Energy_Bin_Pos_88   <= s_Energy_Bin_Pos_88   ;
  o_Energy_Bin_Pos_89   <= s_Energy_Bin_Pos_89   ;
  o_Energy_Bin_Pos_90   <= s_Energy_Bin_Pos_90   ;
  o_Energy_Bin_Pos_91   <= s_Energy_Bin_Pos_91   ;
  o_Energy_Bin_Pos_92   <= s_Energy_Bin_Pos_92   ;
  o_Energy_Bin_Pos_93   <= s_Energy_Bin_Pos_93   ;
  o_Energy_Bin_Pos_94   <= s_Energy_Bin_Pos_94   ;
  o_Energy_Bin_Pos_95   <= s_Energy_Bin_Pos_95   ;
  o_Energy_Bin_Pos_96   <= s_Energy_Bin_Pos_96   ;
  o_Energy_Bin_Pos_97   <= s_Energy_Bin_Pos_97   ;
  o_Energy_Bin_Pos_98   <= s_Energy_Bin_Pos_98   ;
  o_Energy_Bin_Pos_99   <= s_Energy_Bin_Pos_99   ;
  o_Energy_Bin_Pos_100  <= s_Energy_Bin_Pos_100  ;
  o_Energy_Bin_Pos_101  <= s_Energy_Bin_Pos_101  ;
  o_Energy_Bin_Pos_102  <= s_Energy_Bin_Pos_102  ;
  o_Energy_Bin_Pos_103  <= s_Energy_Bin_Pos_103  ;
  o_Energy_Bin_Pos_104  <= s_Energy_Bin_Pos_104  ;
  o_Energy_Bin_Pos_105  <= s_Energy_Bin_Pos_105  ;
  o_Energy_Bin_Pos_106  <= s_Energy_Bin_Pos_106  ;
  o_Energy_Bin_Pos_107  <= s_Energy_Bin_Pos_107  ;
  o_Energy_Bin_Pos_108  <= s_Energy_Bin_Pos_108  ;
  o_Energy_Bin_Pos_109  <= s_Energy_Bin_Pos_109  ;
  o_Energy_Bin_Pos_110  <= s_Energy_Bin_Pos_110  ;
  o_Energy_Bin_Pos_111  <= s_Energy_Bin_Pos_111  ;
  o_Energy_Bin_Pos_112  <= s_Energy_Bin_Pos_112  ;
  o_Energy_Bin_Pos_113  <= s_Energy_Bin_Pos_113  ;
  o_Energy_Bin_Pos_114  <= s_Energy_Bin_Pos_114  ;
  o_Energy_Bin_Pos_115  <= s_Energy_Bin_Pos_115  ;
  o_Energy_Bin_Pos_116  <= s_Energy_Bin_Pos_116  ;
  o_Energy_Bin_Pos_117  <= s_Energy_Bin_Pos_117  ;
  o_Energy_Bin_Pos_118  <= s_Energy_Bin_Pos_118  ;
  o_Energy_Bin_Pos_119  <= s_Energy_Bin_Pos_119  ;
  o_Energy_Bin_Pos_120  <= s_Energy_Bin_Pos_120  ;
  o_Energy_Bin_Pos_121  <= s_Energy_Bin_Pos_121  ;
  o_Energy_Bin_Pos_122  <= s_Energy_Bin_Pos_122  ;
  o_Energy_Bin_Pos_123  <= s_Energy_Bin_Pos_123  ;
  o_Energy_Bin_Pos_124  <= s_Energy_Bin_Pos_124  ;
  o_Energy_Bin_Pos_125  <= s_Energy_Bin_Pos_125  ;
  o_Energy_Bin_Pos_126  <= s_Energy_Bin_Pos_126  ;
  o_Energy_Bin_Pos_127  <= s_Energy_Bin_Pos_127  ;
  o_Energy_Bin_Pos_128  <= s_Energy_Bin_Pos_128  ;
  o_Energy_Bin_Pos_129  <= s_Energy_Bin_Pos_129  ;
  o_Energy_Bin_Pos_130  <= s_Energy_Bin_Pos_130  ;
  o_Energy_Bin_Pos_131  <= s_Energy_Bin_Pos_131  ;
  o_Energy_Bin_Pos_132  <= s_Energy_Bin_Pos_132  ;
  o_Energy_Bin_Pos_133  <= s_Energy_Bin_Pos_133  ;
  o_Energy_Bin_Pos_134  <= s_Energy_Bin_Pos_134  ;
  o_Energy_Bin_Pos_135  <= s_Energy_Bin_Pos_135  ;
  o_Energy_Bin_Pos_136  <= s_Energy_Bin_Pos_136  ;
  o_Energy_Bin_Pos_137  <= s_Energy_Bin_Pos_137  ;
  o_Energy_Bin_Pos_138  <= s_Energy_Bin_Pos_138  ;
  o_Energy_Bin_Pos_139  <= s_Energy_Bin_Pos_139  ;
  o_Energy_Bin_Pos_140  <= s_Energy_Bin_Pos_140  ;
  o_Energy_Bin_Pos_141  <= s_Energy_Bin_Pos_141  ;
  o_Energy_Bin_Pos_142  <= s_Energy_Bin_Pos_142  ;
  o_Energy_Bin_Pos_143  <= s_Energy_Bin_Pos_143  ;
  o_Energy_Bin_Pos_144  <= s_Energy_Bin_Pos_144  ;
  o_Energy_Bin_Pos_145  <= s_Energy_Bin_Pos_145  ;
  o_Energy_Bin_Pos_146  <= s_Energy_Bin_Pos_146  ;
  o_Energy_Bin_Pos_147  <= s_Energy_Bin_Pos_147  ;
  o_Energy_Bin_Pos_148  <= s_Energy_Bin_Pos_148  ;
  o_Energy_Bin_Pos_149  <= s_Energy_Bin_Pos_149  ;
  o_Energy_Bin_Pos_150  <= s_Energy_Bin_Pos_150  ;
  o_Energy_Bin_Pos_151  <= s_Energy_Bin_Pos_151  ;
  o_Energy_Bin_Pos_152  <= s_Energy_Bin_Pos_152  ;
  o_Energy_Bin_Pos_153  <= s_Energy_Bin_Pos_153  ;
  o_Energy_Bin_Pos_154  <= s_Energy_Bin_Pos_154  ;
  o_Energy_Bin_Pos_155  <= s_Energy_Bin_Pos_155  ;
  o_Energy_Bin_Pos_156  <= s_Energy_Bin_Pos_156  ;
  o_Energy_Bin_Pos_157  <= s_Energy_Bin_Pos_157  ;
  o_Energy_Bin_Pos_158  <= s_Energy_Bin_Pos_158  ;
  o_Energy_Bin_Pos_159  <= s_Energy_Bin_Pos_159  ;
  o_Energy_Bin_Pos_160  <= s_Energy_Bin_Pos_160  ;
  o_Energy_Bin_Pos_161  <= s_Energy_Bin_Pos_161  ;
  o_Energy_Bin_Pos_162  <= s_Energy_Bin_Pos_162  ;
  o_Energy_Bin_Pos_163  <= s_Energy_Bin_Pos_163  ;
  o_Energy_Bin_Pos_164  <= s_Energy_Bin_Pos_164  ;
  o_Energy_Bin_Pos_165  <= s_Energy_Bin_Pos_165  ;
  o_Energy_Bin_Pos_166  <= s_Energy_Bin_Pos_166  ;
  o_Energy_Bin_Pos_167  <= s_Energy_Bin_Pos_167  ;
  o_Energy_Bin_Pos_168  <= s_Energy_Bin_Pos_168  ;
  o_Energy_Bin_Pos_169  <= s_Energy_Bin_Pos_169  ;
  o_Energy_Bin_Pos_170  <= s_Energy_Bin_Pos_170  ;
  o_Energy_Bin_Pos_171  <= s_Energy_Bin_Pos_171  ;
  o_Energy_Bin_Pos_172  <= s_Energy_Bin_Pos_172  ;
  o_Energy_Bin_Pos_173  <= s_Energy_Bin_Pos_173  ;
  o_Energy_Bin_Pos_174  <= s_Energy_Bin_Pos_174  ;
  o_Energy_Bin_Pos_175  <= s_Energy_Bin_Pos_175  ;
  o_Energy_Bin_Pos_176  <= s_Energy_Bin_Pos_176  ;
  o_Energy_Bin_Pos_177  <= s_Energy_Bin_Pos_177  ;
  o_Energy_Bin_Pos_178  <= s_Energy_Bin_Pos_178  ;
  o_Energy_Bin_Pos_179  <= s_Energy_Bin_Pos_179  ;
  o_Energy_Bin_Pos_180  <= s_Energy_Bin_Pos_180  ;
  o_Energy_Bin_Pos_181  <= s_Energy_Bin_Pos_181  ;
  o_Energy_Bin_Pos_182  <= s_Energy_Bin_Pos_182  ;
  o_Energy_Bin_Pos_183  <= s_Energy_Bin_Pos_183  ;
  o_Energy_Bin_Pos_184  <= s_Energy_Bin_Pos_184  ;
  o_Energy_Bin_Pos_185  <= s_Energy_Bin_Pos_185  ;
  o_Energy_Bin_Pos_186  <= s_Energy_Bin_Pos_186  ;
  o_Energy_Bin_Pos_187  <= s_Energy_Bin_Pos_187  ;
  o_Energy_Bin_Pos_188  <= s_Energy_Bin_Pos_188  ;
  o_Energy_Bin_Pos_189  <= s_Energy_Bin_Pos_189  ;
  o_Energy_Bin_Pos_190  <= s_Energy_Bin_Pos_190  ;
  o_Energy_Bin_Pos_191  <= s_Energy_Bin_Pos_191  ;
  o_Energy_Bin_Pos_192  <= s_Energy_Bin_Pos_192  ;
  o_Energy_Bin_Pos_193  <= s_Energy_Bin_Pos_193  ;
  o_Energy_Bin_Pos_194  <= s_Energy_Bin_Pos_194  ;
  o_Energy_Bin_Pos_195  <= s_Energy_Bin_Pos_195  ;
  o_Energy_Bin_Pos_196  <= s_Energy_Bin_Pos_196  ;
  o_Energy_Bin_Pos_197  <= s_Energy_Bin_Pos_197  ;
  o_Energy_Bin_Pos_198  <= s_Energy_Bin_Pos_198  ;
  o_Energy_Bin_Pos_199  <= s_Energy_Bin_Pos_199  ;
  o_Energy_Bin_Pos_200  <= s_Energy_Bin_Pos_200  ;
  o_Energy_Bin_Pos_201  <= s_Energy_Bin_Pos_201  ;
  o_Energy_Bin_Pos_202  <= s_Energy_Bin_Pos_202  ;
  o_Energy_Bin_Pos_203  <= s_Energy_Bin_Pos_203  ;
  o_Energy_Bin_Pos_204  <= s_Energy_Bin_Pos_204  ;
  o_Energy_Bin_Pos_205  <= s_Energy_Bin_Pos_205  ;
  o_Energy_Bin_Pos_206  <= s_Energy_Bin_Pos_206  ;
  o_Energy_Bin_Pos_207  <= s_Energy_Bin_Pos_207  ;
  o_Energy_Bin_Pos_208  <= s_Energy_Bin_Pos_208  ;
  o_Energy_Bin_Pos_209  <= s_Energy_Bin_Pos_209  ;
  o_Energy_Bin_Pos_210  <= s_Energy_Bin_Pos_210  ;
  o_Energy_Bin_Pos_211  <= s_Energy_Bin_Pos_211  ;
  o_Energy_Bin_Pos_212  <= s_Energy_Bin_Pos_212  ;
  o_Energy_Bin_Pos_213  <= s_Energy_Bin_Pos_213  ;
  o_Energy_Bin_Pos_214  <= s_Energy_Bin_Pos_214  ;
  o_Energy_Bin_Pos_215  <= s_Energy_Bin_Pos_215  ;
  o_Energy_Bin_Pos_216  <= s_Energy_Bin_Pos_216  ;
  o_Energy_Bin_Pos_217  <= s_Energy_Bin_Pos_217  ;
  o_Energy_Bin_Pos_218  <= s_Energy_Bin_Pos_218  ;
  o_Energy_Bin_Pos_219  <= s_Energy_Bin_Pos_219  ;
  o_Energy_Bin_Pos_220  <= s_Energy_Bin_Pos_220  ;
  o_Energy_Bin_Pos_221  <= s_Energy_Bin_Pos_221  ;
  o_Energy_Bin_Pos_222  <= s_Energy_Bin_Pos_222  ;
  o_Energy_Bin_Pos_223  <= s_Energy_Bin_Pos_223  ;
  o_Energy_Bin_Pos_224  <= s_Energy_Bin_Pos_224  ;
  o_Energy_Bin_Pos_225  <= s_Energy_Bin_Pos_225  ;
  o_Energy_Bin_Pos_226  <= s_Energy_Bin_Pos_226  ;
  o_Energy_Bin_Pos_227  <= s_Energy_Bin_Pos_227  ;
  o_Energy_Bin_Pos_228  <= s_Energy_Bin_Pos_228  ;
  o_Energy_Bin_Pos_229  <= s_Energy_Bin_Pos_229  ;
  o_Energy_Bin_Pos_230  <= s_Energy_Bin_Pos_230  ;
  o_Energy_Bin_Pos_231  <= s_Energy_Bin_Pos_231  ;
  o_Energy_Bin_Pos_232  <= s_Energy_Bin_Pos_232  ;
  o_Energy_Bin_Pos_233  <= s_Energy_Bin_Pos_233  ;
  o_Energy_Bin_Pos_234  <= s_Energy_Bin_Pos_234  ;
  o_Energy_Bin_Pos_235  <= s_Energy_Bin_Pos_235  ;
  o_Energy_Bin_Pos_236  <= s_Energy_Bin_Pos_236  ;
  o_Energy_Bin_Pos_237  <= s_Energy_Bin_Pos_237  ;
  o_Energy_Bin_Pos_238  <= s_Energy_Bin_Pos_238  ;
  o_Energy_Bin_Pos_239  <= s_Energy_Bin_Pos_239  ;
  o_Energy_Bin_Pos_240  <= s_Energy_Bin_Pos_240  ;
  o_Energy_Bin_Pos_241  <= s_Energy_Bin_Pos_241  ;
  o_Energy_Bin_Pos_242  <= s_Energy_Bin_Pos_242  ;
  o_Energy_Bin_Pos_243  <= s_Energy_Bin_Pos_243  ;
  o_Energy_Bin_Pos_244  <= s_Energy_Bin_Pos_244  ;
  o_Energy_Bin_Pos_245  <= s_Energy_Bin_Pos_245  ;
  o_Energy_Bin_Pos_246  <= s_Energy_Bin_Pos_246  ;
  o_Energy_Bin_Pos_247  <= s_Energy_Bin_Pos_247  ;
  o_Energy_Bin_Pos_248  <= s_Energy_Bin_Pos_248  ;
  o_Energy_Bin_Pos_249  <= s_Energy_Bin_Pos_249  ;
  o_Energy_Bin_Pos_250  <= s_Energy_Bin_Pos_250  ;
  o_Energy_Bin_Pos_251  <= s_Energy_Bin_Pos_251  ;
  o_Energy_Bin_Pos_252  <= s_Energy_Bin_Pos_252  ;
  o_Energy_Bin_Pos_253  <= s_Energy_Bin_Pos_253  ;
  o_Energy_Bin_Pos_254  <= s_Energy_Bin_Pos_254  ;
  o_Energy_Bin_Pos_255  <= s_Energy_Bin_Pos_255  ;
  o_Energy_Bin_Pos_256  <= s_Energy_Bin_Pos_256  ;
  o_Energy_Bin_Pos_257  <= s_Energy_Bin_Pos_257  ;
  o_Energy_Bin_Pos_258  <= s_Energy_Bin_Pos_258  ;
  o_Energy_Bin_Pos_259  <= s_Energy_Bin_Pos_259  ;
  o_Energy_Bin_Pos_260  <= s_Energy_Bin_Pos_260  ;
  o_Energy_Bin_Pos_261  <= s_Energy_Bin_Pos_261  ;
  o_Energy_Bin_Pos_262  <= s_Energy_Bin_Pos_262  ;
  o_Energy_Bin_Pos_263  <= s_Energy_Bin_Pos_263  ;
  o_Energy_Bin_Pos_264  <= s_Energy_Bin_Pos_264  ;
  o_Energy_Bin_Pos_265  <= s_Energy_Bin_Pos_265  ;
  o_Energy_Bin_Pos_266  <= s_Energy_Bin_Pos_266  ;
  o_Energy_Bin_Pos_267  <= s_Energy_Bin_Pos_267  ;
  o_Energy_Bin_Pos_268  <= s_Energy_Bin_Pos_268  ;
  o_Energy_Bin_Pos_269  <= s_Energy_Bin_Pos_269  ;
  o_Energy_Bin_Pos_270  <= s_Energy_Bin_Pos_270  ;
  o_Energy_Bin_Pos_271  <= s_Energy_Bin_Pos_271  ;
  o_Energy_Bin_Pos_272  <= s_Energy_Bin_Pos_272  ;
  o_Energy_Bin_Pos_273  <= s_Energy_Bin_Pos_273  ;
  o_Energy_Bin_Pos_274  <= s_Energy_Bin_Pos_274  ;
  o_Energy_Bin_Pos_275  <= s_Energy_Bin_Pos_275  ;
  o_Energy_Bin_Pos_276  <= s_Energy_Bin_Pos_276  ;
  o_Energy_Bin_Pos_277  <= s_Energy_Bin_Pos_277  ;
  o_Energy_Bin_Pos_278  <= s_Energy_Bin_Pos_278  ;
  o_Energy_Bin_Pos_279  <= s_Energy_Bin_Pos_279  ;
  o_Energy_Bin_Pos_280  <= s_Energy_Bin_Pos_280  ;
  o_Energy_Bin_Pos_281  <= s_Energy_Bin_Pos_281  ;
  o_Energy_Bin_Pos_282  <= s_Energy_Bin_Pos_282  ;
  o_Energy_Bin_Pos_283  <= s_Energy_Bin_Pos_283  ;
  o_Energy_Bin_Pos_284  <= s_Energy_Bin_Pos_284  ;
  o_Energy_Bin_Pos_285  <= s_Energy_Bin_Pos_285  ;
  o_Energy_Bin_Pos_286  <= s_Energy_Bin_Pos_286  ;
  o_Energy_Bin_Pos_287  <= s_Energy_Bin_Pos_287  ;
  o_Energy_Bin_Pos_288  <= s_Energy_Bin_Pos_288  ;
  o_Energy_Bin_Pos_289  <= s_Energy_Bin_Pos_289  ;
  o_Energy_Bin_Pos_290  <= s_Energy_Bin_Pos_290  ;
  o_Energy_Bin_Pos_291  <= s_Energy_Bin_Pos_291  ;
  o_Energy_Bin_Pos_292  <= s_Energy_Bin_Pos_292  ;
  o_Energy_Bin_Pos_293  <= s_Energy_Bin_Pos_293  ;
  o_Energy_Bin_Pos_294  <= s_Energy_Bin_Pos_294  ;
  o_Energy_Bin_Pos_295  <= s_Energy_Bin_Pos_295  ;
  o_Energy_Bin_Pos_296  <= s_Energy_Bin_Pos_296  ;
  o_Energy_Bin_Pos_297  <= s_Energy_Bin_Pos_297  ;
  o_Energy_Bin_Pos_298  <= s_Energy_Bin_Pos_298  ;
  o_Energy_Bin_Pos_299  <= s_Energy_Bin_Pos_299  ;
  o_Energy_Bin_Pos_300  <= s_Energy_Bin_Pos_300  ;
  o_Energy_Bin_Pos_301  <= s_Energy_Bin_Pos_301  ;
  o_Energy_Bin_Pos_302  <= s_Energy_Bin_Pos_302  ;
  o_Energy_Bin_Pos_303  <= s_Energy_Bin_Pos_303  ;
  o_Energy_Bin_Pos_304  <= s_Energy_Bin_Pos_304  ;
  o_Energy_Bin_Pos_305  <= s_Energy_Bin_Pos_305  ;
  o_Energy_Bin_Pos_306  <= s_Energy_Bin_Pos_306  ;
  o_Energy_Bin_Pos_307  <= s_Energy_Bin_Pos_307  ;
  o_Energy_Bin_Pos_308  <= s_Energy_Bin_Pos_308  ;
  o_Energy_Bin_Pos_309  <= s_Energy_Bin_Pos_309  ;
  o_Energy_Bin_Pos_310  <= s_Energy_Bin_Pos_310  ;
  o_Energy_Bin_Pos_311  <= s_Energy_Bin_Pos_311  ;
  o_Energy_Bin_Pos_312  <= s_Energy_Bin_Pos_312  ;
  o_Energy_Bin_Pos_313  <= s_Energy_Bin_Pos_313  ;
  o_Energy_Bin_Pos_314  <= s_Energy_Bin_Pos_314  ;
  o_Energy_Bin_Pos_315  <= s_Energy_Bin_Pos_315  ;
  o_Energy_Bin_Pos_316  <= s_Energy_Bin_Pos_316  ;
  o_Energy_Bin_Pos_317  <= s_Energy_Bin_Pos_317  ;
  o_Energy_Bin_Pos_318  <= s_Energy_Bin_Pos_318  ;
  o_Energy_Bin_Pos_319  <= s_Energy_Bin_Pos_319  ;
  o_Energy_Bin_Pos_320  <= s_Energy_Bin_Pos_320  ;
  o_Energy_Bin_Pos_321  <= s_Energy_Bin_Pos_321  ;
  o_Energy_Bin_Pos_322  <= s_Energy_Bin_Pos_322  ;
  o_Energy_Bin_Pos_323  <= s_Energy_Bin_Pos_323  ;
  o_Energy_Bin_Pos_324  <= s_Energy_Bin_Pos_324  ;
  o_Energy_Bin_Pos_325  <= s_Energy_Bin_Pos_325  ;
  o_Energy_Bin_Pos_326  <= s_Energy_Bin_Pos_326  ;
  o_Energy_Bin_Pos_327  <= s_Energy_Bin_Pos_327  ;
  o_Energy_Bin_Pos_328  <= s_Energy_Bin_Pos_328  ;
  o_Energy_Bin_Pos_329  <= s_Energy_Bin_Pos_329  ;
  o_Energy_Bin_Pos_330  <= s_Energy_Bin_Pos_330  ;
  o_Energy_Bin_Pos_331  <= s_Energy_Bin_Pos_331  ;
  o_Energy_Bin_Pos_332  <= s_Energy_Bin_Pos_332  ;
  o_Energy_Bin_Pos_333  <= s_Energy_Bin_Pos_333  ;
  o_Energy_Bin_Pos_334  <= s_Energy_Bin_Pos_334  ;
  o_Energy_Bin_Pos_335  <= s_Energy_Bin_Pos_335  ;
  o_Energy_Bin_Pos_336  <= s_Energy_Bin_Pos_336  ;
  o_Energy_Bin_Pos_337  <= s_Energy_Bin_Pos_337  ;
  o_Energy_Bin_Pos_338  <= s_Energy_Bin_Pos_338  ;
  o_Energy_Bin_Pos_339  <= s_Energy_Bin_Pos_339  ;
  o_Energy_Bin_Pos_340  <= s_Energy_Bin_Pos_340  ;
  o_Energy_Bin_Pos_341  <= s_Energy_Bin_Pos_341  ;
  o_Energy_Bin_Pos_342  <= s_Energy_Bin_Pos_342  ;
  o_Energy_Bin_Pos_343  <= s_Energy_Bin_Pos_343  ;
  o_Energy_Bin_Pos_344  <= s_Energy_Bin_Pos_344  ;
  o_Energy_Bin_Pos_345  <= s_Energy_Bin_Pos_345  ;
  o_Energy_Bin_Pos_346  <= s_Energy_Bin_Pos_346  ;
  o_Energy_Bin_Pos_347  <= s_Energy_Bin_Pos_347  ;
  o_Energy_Bin_Pos_348  <= s_Energy_Bin_Pos_348  ;
  o_Energy_Bin_Pos_349  <= s_Energy_Bin_Pos_349  ;
  o_Energy_Bin_Pos_350  <= s_Energy_Bin_Pos_350  ;
  o_Energy_Bin_Pos_351  <= s_Energy_Bin_Pos_351  ;
  o_Energy_Bin_Pos_352  <= s_Energy_Bin_Pos_352  ;
  o_Energy_Bin_Pos_353  <= s_Energy_Bin_Pos_353  ;
  o_Energy_Bin_Pos_354  <= s_Energy_Bin_Pos_354  ;
  o_Energy_Bin_Pos_355  <= s_Energy_Bin_Pos_355  ;
  o_Energy_Bin_Pos_356  <= s_Energy_Bin_Pos_356  ;
  o_Energy_Bin_Pos_357  <= s_Energy_Bin_Pos_357  ;
  o_Energy_Bin_Pos_358  <= s_Energy_Bin_Pos_358  ;
  o_Energy_Bin_Pos_359  <= s_Energy_Bin_Pos_359  ;
  o_Energy_Bin_Pos_360  <= s_Energy_Bin_Pos_360  ;
  o_Energy_Bin_Pos_361  <= s_Energy_Bin_Pos_361  ;
  o_Energy_Bin_Pos_362  <= s_Energy_Bin_Pos_362  ;
  o_Energy_Bin_Pos_363  <= s_Energy_Bin_Pos_363  ;
  o_Energy_Bin_Pos_364  <= s_Energy_Bin_Pos_364  ;
  o_Energy_Bin_Pos_365  <= s_Energy_Bin_Pos_365  ;
  o_Energy_Bin_Pos_366  <= s_Energy_Bin_Pos_366  ;
  o_Energy_Bin_Pos_367  <= s_Energy_Bin_Pos_367  ;
  o_Energy_Bin_Pos_368  <= s_Energy_Bin_Pos_368  ;
  o_Energy_Bin_Pos_369  <= s_Energy_Bin_Pos_369  ;
  o_Energy_Bin_Pos_370  <= s_Energy_Bin_Pos_370  ;
  o_Energy_Bin_Pos_371  <= s_Energy_Bin_Pos_371  ;
  o_Energy_Bin_Pos_372  <= s_Energy_Bin_Pos_372  ;
  o_Energy_Bin_Pos_373  <= s_Energy_Bin_Pos_373  ;
  o_Energy_Bin_Pos_374  <= s_Energy_Bin_Pos_374  ;
  o_Energy_Bin_Pos_375  <= s_Energy_Bin_Pos_375  ;
  o_Energy_Bin_Pos_376  <= s_Energy_Bin_Pos_376  ;
  o_Energy_Bin_Pos_377  <= s_Energy_Bin_Pos_377  ;
  o_Energy_Bin_Pos_378  <= s_Energy_Bin_Pos_378  ;
  o_Energy_Bin_Pos_379  <= s_Energy_Bin_Pos_379  ;
  o_Energy_Bin_Pos_380  <= s_Energy_Bin_Pos_380  ;
  o_Energy_Bin_Pos_381  <= s_Energy_Bin_Pos_381  ;
  o_Energy_Bin_Pos_382  <= s_Energy_Bin_Pos_382  ;
  o_Energy_Bin_Pos_383  <= s_Energy_Bin_Pos_383  ;
  o_Energy_Bin_Pos_384  <= s_Energy_Bin_Pos_384  ;
  o_Energy_Bin_Pos_385  <= s_Energy_Bin_Pos_385  ;
  o_Energy_Bin_Pos_386  <= s_Energy_Bin_Pos_386  ;
  o_Energy_Bin_Pos_387  <= s_Energy_Bin_Pos_387  ;
  o_Energy_Bin_Pos_388  <= s_Energy_Bin_Pos_388  ;
  o_Energy_Bin_Pos_389  <= s_Energy_Bin_Pos_389  ;
  o_Energy_Bin_Pos_390  <= s_Energy_Bin_Pos_390  ;
  o_Energy_Bin_Pos_391  <= s_Energy_Bin_Pos_391  ;
  o_Energy_Bin_Pos_392  <= s_Energy_Bin_Pos_392  ;
  o_Energy_Bin_Pos_393  <= s_Energy_Bin_Pos_393  ;
  o_Energy_Bin_Pos_394  <= s_Energy_Bin_Pos_394  ;
  o_Energy_Bin_Pos_395  <= s_Energy_Bin_Pos_395  ;
  o_Energy_Bin_Pos_396  <= s_Energy_Bin_Pos_396  ;
  o_Energy_Bin_Pos_397  <= s_Energy_Bin_Pos_397  ;
  o_Energy_Bin_Pos_398  <= s_Energy_Bin_Pos_398  ;
  o_Energy_Bin_Pos_399  <= s_Energy_Bin_Pos_399  ;
  o_Energy_Bin_Pos_400  <= s_Energy_Bin_Pos_400  ;
  o_Energy_Bin_Pos_401  <= s_Energy_Bin_Pos_401  ;
  o_Energy_Bin_Pos_402  <= s_Energy_Bin_Pos_402  ;
  o_Energy_Bin_Pos_403  <= s_Energy_Bin_Pos_403  ;
  o_Energy_Bin_Pos_404  <= s_Energy_Bin_Pos_404  ;
  o_Energy_Bin_Pos_405  <= s_Energy_Bin_Pos_405  ;
  o_Energy_Bin_Pos_406  <= s_Energy_Bin_Pos_406  ;
  o_Energy_Bin_Pos_407  <= s_Energy_Bin_Pos_407  ;
  o_Energy_Bin_Pos_408  <= s_Energy_Bin_Pos_408  ;
  o_Energy_Bin_Pos_409  <= s_Energy_Bin_Pos_409  ;
  o_Energy_Bin_Pos_410  <= s_Energy_Bin_Pos_410  ;
  o_Energy_Bin_Pos_411  <= s_Energy_Bin_Pos_411  ;
  o_Energy_Bin_Pos_412  <= s_Energy_Bin_Pos_412  ;
  o_Energy_Bin_Pos_413  <= s_Energy_Bin_Pos_413  ;
  o_Energy_Bin_Pos_414  <= s_Energy_Bin_Pos_414  ;
  o_Energy_Bin_Pos_415  <= s_Energy_Bin_Pos_415  ;
  o_Energy_Bin_Pos_416  <= s_Energy_Bin_Pos_416  ;
  o_Energy_Bin_Pos_417  <= s_Energy_Bin_Pos_417  ;
  o_Energy_Bin_Pos_418  <= s_Energy_Bin_Pos_418  ;
  o_Energy_Bin_Pos_419  <= s_Energy_Bin_Pos_419  ;
  o_Energy_Bin_Pos_420  <= s_Energy_Bin_Pos_420  ;
  o_Energy_Bin_Pos_421  <= s_Energy_Bin_Pos_421  ;
  o_Energy_Bin_Pos_422  <= s_Energy_Bin_Pos_422  ;
  o_Energy_Bin_Pos_423  <= s_Energy_Bin_Pos_423  ;
  o_Energy_Bin_Pos_424  <= s_Energy_Bin_Pos_424  ;
  o_Energy_Bin_Pos_425  <= s_Energy_Bin_Pos_425  ;
  o_Energy_Bin_Pos_426  <= s_Energy_Bin_Pos_426  ;
  o_Energy_Bin_Pos_427  <= s_Energy_Bin_Pos_427  ;
  o_Energy_Bin_Pos_428  <= s_Energy_Bin_Pos_428  ;
  o_Energy_Bin_Pos_429  <= s_Energy_Bin_Pos_429  ;
  o_Energy_Bin_Pos_430  <= s_Energy_Bin_Pos_430  ;
  o_Energy_Bin_Pos_431  <= s_Energy_Bin_Pos_431  ;
  o_Energy_Bin_Pos_432  <= s_Energy_Bin_Pos_432  ;
  o_Energy_Bin_Pos_433  <= s_Energy_Bin_Pos_433  ;
  o_Energy_Bin_Pos_434  <= s_Energy_Bin_Pos_434  ;
  o_Energy_Bin_Pos_435  <= s_Energy_Bin_Pos_435  ;
  o_Energy_Bin_Pos_436  <= s_Energy_Bin_Pos_436  ;
  o_Energy_Bin_Pos_437  <= s_Energy_Bin_Pos_437  ;
  o_Energy_Bin_Pos_438  <= s_Energy_Bin_Pos_438  ;
  o_Energy_Bin_Pos_439  <= s_Energy_Bin_Pos_439  ;
  o_Energy_Bin_Pos_440  <= s_Energy_Bin_Pos_440  ;
  o_Energy_Bin_Pos_441  <= s_Energy_Bin_Pos_441  ;
  o_Energy_Bin_Pos_442  <= s_Energy_Bin_Pos_442  ;
  o_Energy_Bin_Pos_443  <= s_Energy_Bin_Pos_443  ;
  o_Energy_Bin_Pos_444  <= s_Energy_Bin_Pos_444  ;
  o_Energy_Bin_Pos_445  <= s_Energy_Bin_Pos_445  ;
  o_Energy_Bin_Pos_446  <= s_Energy_Bin_Pos_446  ;
  o_Energy_Bin_Pos_447  <= s_Energy_Bin_Pos_447  ;
  o_Energy_Bin_Pos_448  <= s_Energy_Bin_Pos_448  ;
  o_Energy_Bin_Pos_449  <= s_Energy_Bin_Pos_449  ;
  o_Energy_Bin_Pos_450  <= s_Energy_Bin_Pos_450  ;
  o_Energy_Bin_Pos_451  <= s_Energy_Bin_Pos_451  ;
  o_Energy_Bin_Pos_452  <= s_Energy_Bin_Pos_452  ;
  o_Energy_Bin_Pos_453  <= s_Energy_Bin_Pos_453  ;
  o_Energy_Bin_Pos_454  <= s_Energy_Bin_Pos_454  ;
  o_Energy_Bin_Pos_455  <= s_Energy_Bin_Pos_455  ;
  o_Energy_Bin_Pos_456  <= s_Energy_Bin_Pos_456  ;
  o_Energy_Bin_Pos_457  <= s_Energy_Bin_Pos_457  ;
  o_Energy_Bin_Pos_458  <= s_Energy_Bin_Pos_458  ;
  o_Energy_Bin_Pos_459  <= s_Energy_Bin_Pos_459  ;
  o_Energy_Bin_Pos_460  <= s_Energy_Bin_Pos_460  ;
  o_Energy_Bin_Pos_461  <= s_Energy_Bin_Pos_461  ;
  o_Energy_Bin_Pos_462  <= s_Energy_Bin_Pos_462  ;
  o_Energy_Bin_Pos_463  <= s_Energy_Bin_Pos_463  ;
  o_Energy_Bin_Pos_464  <= s_Energy_Bin_Pos_464  ;
  o_Energy_Bin_Pos_465  <= s_Energy_Bin_Pos_465  ;
  o_Energy_Bin_Pos_466  <= s_Energy_Bin_Pos_466  ;
  o_Energy_Bin_Pos_467  <= s_Energy_Bin_Pos_467  ;
  o_Energy_Bin_Pos_468  <= s_Energy_Bin_Pos_468  ;
  o_Energy_Bin_Pos_469  <= s_Energy_Bin_Pos_469  ;
  o_Energy_Bin_Pos_470  <= s_Energy_Bin_Pos_470  ;
  o_Energy_Bin_Pos_471  <= s_Energy_Bin_Pos_471  ;
  o_Energy_Bin_Pos_472  <= s_Energy_Bin_Pos_472  ;
  o_Energy_Bin_Pos_473  <= s_Energy_Bin_Pos_473  ;
  o_Energy_Bin_Pos_474  <= s_Energy_Bin_Pos_474  ;
  o_Energy_Bin_Pos_475  <= s_Energy_Bin_Pos_475  ;
  o_Energy_Bin_Pos_476  <= s_Energy_Bin_Pos_476  ;
  o_Energy_Bin_Pos_477  <= s_Energy_Bin_Pos_477  ;
  o_Energy_Bin_Pos_478  <= s_Energy_Bin_Pos_478  ;
  o_Energy_Bin_Pos_479  <= s_Energy_Bin_Pos_479  ;
  o_Energy_Bin_Pos_480  <= s_Energy_Bin_Pos_480  ;
  o_Energy_Bin_Pos_481  <= s_Energy_Bin_Pos_481  ;
  o_Energy_Bin_Pos_482  <= s_Energy_Bin_Pos_482  ;
  o_Energy_Bin_Pos_483  <= s_Energy_Bin_Pos_483  ;
  o_Energy_Bin_Pos_484  <= s_Energy_Bin_Pos_484  ;
  o_Energy_Bin_Pos_485  <= s_Energy_Bin_Pos_485  ;
  o_Energy_Bin_Pos_486  <= s_Energy_Bin_Pos_486  ;
  o_Energy_Bin_Pos_487  <= s_Energy_Bin_Pos_487  ;
  o_Energy_Bin_Pos_488  <= s_Energy_Bin_Pos_488  ;
  o_Energy_Bin_Pos_489  <= s_Energy_Bin_Pos_489  ;
  o_Energy_Bin_Pos_490  <= s_Energy_Bin_Pos_490  ;
  o_Energy_Bin_Pos_491  <= s_Energy_Bin_Pos_491  ;
  o_Energy_Bin_Pos_492  <= s_Energy_Bin_Pos_492  ;
  o_Energy_Bin_Pos_493  <= s_Energy_Bin_Pos_493  ;
  o_Energy_Bin_Pos_494  <= s_Energy_Bin_Pos_494  ;
  o_Energy_Bin_Pos_495  <= s_Energy_Bin_Pos_495  ;
  o_Energy_Bin_Pos_496  <= s_Energy_Bin_Pos_496  ;
  o_Energy_Bin_Pos_497  <= s_Energy_Bin_Pos_497  ;
  o_Energy_Bin_Pos_498  <= s_Energy_Bin_Pos_498  ;
  o_Energy_Bin_Pos_499  <= s_Energy_Bin_Pos_499  ;
  o_Energy_Bin_Pos_500  <= s_Energy_Bin_Pos_500  ;
  o_Energy_Bin_Pos_501  <= s_Energy_Bin_Pos_501  ;
  o_Energy_Bin_Pos_502  <= s_Energy_Bin_Pos_502  ;
  o_Energy_Bin_Pos_503  <= s_Energy_Bin_Pos_503  ;
  o_Energy_Bin_Pos_504  <= s_Energy_Bin_Pos_504  ;
  o_Energy_Bin_Pos_505  <= s_Energy_Bin_Pos_505  ;
  o_Energy_Bin_Pos_506  <= s_Energy_Bin_Pos_506  ;
  o_Energy_Bin_Pos_507  <= s_Energy_Bin_Pos_507  ;
  o_Energy_Bin_Pos_508  <= s_Energy_Bin_Pos_508  ;
  o_Energy_Bin_Pos_509  <= s_Energy_Bin_Pos_509  ;
  o_Energy_Bin_Pos_510  <= s_Energy_Bin_Pos_510  ;
  o_Energy_Bin_Pos_511  <= s_Energy_Bin_Pos_511  ;
  o_Energy_Bin_Pos_512  <= s_Energy_Bin_Pos_512  ;
  o_Energy_Bin_Pos_513  <= s_Energy_Bin_Pos_513  ;
  o_Energy_Bin_Pos_514  <= s_Energy_Bin_Pos_514  ;
  o_Energy_Bin_Pos_515  <= s_Energy_Bin_Pos_515  ;
  o_Energy_Bin_Pos_516  <= s_Energy_Bin_Pos_516  ;
  o_Energy_Bin_Pos_517  <= s_Energy_Bin_Pos_517  ;
  o_Energy_Bin_Pos_518  <= s_Energy_Bin_Pos_518  ;
  o_Energy_Bin_Pos_519  <= s_Energy_Bin_Pos_519  ;
  o_Energy_Bin_Pos_520  <= s_Energy_Bin_Pos_520  ;
  o_Energy_Bin_Pos_521  <= s_Energy_Bin_Pos_521  ;
  o_Energy_Bin_Pos_522  <= s_Energy_Bin_Pos_522  ;
  o_Energy_Bin_Pos_523  <= s_Energy_Bin_Pos_523  ;
  o_Energy_Bin_Pos_524  <= s_Energy_Bin_Pos_524  ;
  o_Energy_Bin_Pos_525  <= s_Energy_Bin_Pos_525  ;
  o_Energy_Bin_Pos_526  <= s_Energy_Bin_Pos_526  ;
  o_Energy_Bin_Pos_527  <= s_Energy_Bin_Pos_527  ;
  o_Energy_Bin_Pos_528  <= s_Energy_Bin_Pos_528  ;
  o_Energy_Bin_Pos_529  <= s_Energy_Bin_Pos_529  ;
  o_Energy_Bin_Pos_530  <= s_Energy_Bin_Pos_530  ;
  o_Energy_Bin_Pos_531  <= s_Energy_Bin_Pos_531  ;
  o_Energy_Bin_Pos_532  <= s_Energy_Bin_Pos_532  ;
  o_Energy_Bin_Pos_533  <= s_Energy_Bin_Pos_533  ;
  o_Energy_Bin_Pos_534  <= s_Energy_Bin_Pos_534  ;
  o_Energy_Bin_Pos_535  <= s_Energy_Bin_Pos_535  ;
  o_Energy_Bin_Pos_536  <= s_Energy_Bin_Pos_536  ;
  o_Energy_Bin_Pos_537  <= s_Energy_Bin_Pos_537  ;
  o_Energy_Bin_Pos_538  <= s_Energy_Bin_Pos_538  ;
  o_Energy_Bin_Pos_539  <= s_Energy_Bin_Pos_539  ;
  o_Energy_Bin_Pos_540  <= s_Energy_Bin_Pos_540  ;
  o_Energy_Bin_Pos_541  <= s_Energy_Bin_Pos_541  ;
  o_Energy_Bin_Pos_542  <= s_Energy_Bin_Pos_542  ;
  o_Energy_Bin_Pos_543  <= s_Energy_Bin_Pos_543  ;
  o_Energy_Bin_Pos_544  <= s_Energy_Bin_Pos_544  ;
  o_Energy_Bin_Pos_545  <= s_Energy_Bin_Pos_545  ;
  o_Energy_Bin_Pos_546  <= s_Energy_Bin_Pos_546  ;
  o_Energy_Bin_Pos_547  <= s_Energy_Bin_Pos_547  ;
  o_Energy_Bin_Pos_548  <= s_Energy_Bin_Pos_548  ;
  o_Energy_Bin_Pos_549  <= s_Energy_Bin_Pos_549  ;
  o_Energy_Bin_Pos_550  <= s_Energy_Bin_Pos_550  ;
  o_Energy_Bin_Pos_551  <= s_Energy_Bin_Pos_551  ;
  o_Energy_Bin_Pos_552  <= s_Energy_Bin_Pos_552  ;
  o_Energy_Bin_Pos_553  <= s_Energy_Bin_Pos_553  ;
  o_Energy_Bin_Pos_554  <= s_Energy_Bin_Pos_554  ;
  o_Energy_Bin_Pos_555  <= s_Energy_Bin_Pos_555  ;
  o_Energy_Bin_Pos_556  <= s_Energy_Bin_Pos_556  ;
  o_Energy_Bin_Pos_557  <= s_Energy_Bin_Pos_557  ;
  o_Energy_Bin_Pos_558  <= s_Energy_Bin_Pos_558  ;
  o_Energy_Bin_Pos_559  <= s_Energy_Bin_Pos_559  ;
  o_Energy_Bin_Pos_560  <= s_Energy_Bin_Pos_560  ;
  o_Energy_Bin_Pos_561  <= s_Energy_Bin_Pos_561  ;
  o_Energy_Bin_Pos_562  <= s_Energy_Bin_Pos_562  ;
  o_Energy_Bin_Pos_563  <= s_Energy_Bin_Pos_563  ;
  o_Energy_Bin_Pos_564  <= s_Energy_Bin_Pos_564  ;
  o_Energy_Bin_Pos_565  <= s_Energy_Bin_Pos_565  ;
  o_Energy_Bin_Pos_566  <= s_Energy_Bin_Pos_566  ;
  o_Energy_Bin_Pos_567  <= s_Energy_Bin_Pos_567  ;
  o_Energy_Bin_Pos_568  <= s_Energy_Bin_Pos_568  ;
  o_Energy_Bin_Pos_569  <= s_Energy_Bin_Pos_569  ;
  o_Energy_Bin_Pos_570  <= s_Energy_Bin_Pos_570  ;
  o_Energy_Bin_Pos_571  <= s_Energy_Bin_Pos_571  ;
  o_Energy_Bin_Pos_572  <= s_Energy_Bin_Pos_572  ;
  o_Energy_Bin_Pos_573  <= s_Energy_Bin_Pos_573  ;
  o_Energy_Bin_Pos_574  <= s_Energy_Bin_Pos_574  ;
  o_Energy_Bin_Pos_575  <= s_Energy_Bin_Pos_575  ;
  o_Energy_Bin_Pos_576  <= s_Energy_Bin_Pos_576  ;
  o_Energy_Bin_Pos_577  <= s_Energy_Bin_Pos_577  ;
  o_Energy_Bin_Pos_578  <= s_Energy_Bin_Pos_578  ;
  o_Energy_Bin_Pos_579  <= s_Energy_Bin_Pos_579  ;
  o_Energy_Bin_Pos_580  <= s_Energy_Bin_Pos_580  ;
  o_Energy_Bin_Pos_581  <= s_Energy_Bin_Pos_581  ;
  o_Energy_Bin_Pos_582  <= s_Energy_Bin_Pos_582  ;
  o_Energy_Bin_Pos_583  <= s_Energy_Bin_Pos_583  ;
  o_Energy_Bin_Pos_584  <= s_Energy_Bin_Pos_584  ;
  o_Energy_Bin_Pos_585  <= s_Energy_Bin_Pos_585  ;
  o_Energy_Bin_Pos_586  <= s_Energy_Bin_Pos_586  ;
  o_Energy_Bin_Pos_587  <= s_Energy_Bin_Pos_587  ;
  o_Energy_Bin_Pos_588  <= s_Energy_Bin_Pos_588  ;
  o_Energy_Bin_Pos_589  <= s_Energy_Bin_Pos_589  ;
  o_Energy_Bin_Pos_590  <= s_Energy_Bin_Pos_590  ;
  o_Energy_Bin_Pos_591  <= s_Energy_Bin_Pos_591  ;
  o_Energy_Bin_Pos_592  <= s_Energy_Bin_Pos_592  ;
  o_Energy_Bin_Pos_593  <= s_Energy_Bin_Pos_593  ;
  o_Energy_Bin_Pos_594  <= s_Energy_Bin_Pos_594  ;
  o_Energy_Bin_Pos_595  <= s_Energy_Bin_Pos_595  ;
  o_Energy_Bin_Pos_596  <= s_Energy_Bin_Pos_596  ;
  o_Energy_Bin_Pos_597  <= s_Energy_Bin_Pos_597  ;
  o_Energy_Bin_Pos_598  <= s_Energy_Bin_Pos_598  ;
  o_Energy_Bin_Pos_599  <= s_Energy_Bin_Pos_599  ;
  o_Energy_Bin_Pos_600  <= s_Energy_Bin_Pos_600  ;
  o_Energy_Bin_Pos_601  <= s_Energy_Bin_Pos_601  ;
  o_Energy_Bin_Pos_602  <= s_Energy_Bin_Pos_602  ;
  o_Energy_Bin_Pos_603  <= s_Energy_Bin_Pos_603  ;
  o_Energy_Bin_Pos_604  <= s_Energy_Bin_Pos_604  ;
  o_Energy_Bin_Pos_605  <= s_Energy_Bin_Pos_605  ;
  o_Energy_Bin_Pos_606  <= s_Energy_Bin_Pos_606  ;
  o_Energy_Bin_Pos_607  <= s_Energy_Bin_Pos_607  ;
  o_Energy_Bin_Pos_608  <= s_Energy_Bin_Pos_608  ;
  o_Energy_Bin_Pos_609  <= s_Energy_Bin_Pos_609  ;
  o_Energy_Bin_Pos_610  <= s_Energy_Bin_Pos_610  ;
  o_Energy_Bin_Pos_611  <= s_Energy_Bin_Pos_611  ;
  o_Energy_Bin_Pos_612  <= s_Energy_Bin_Pos_612  ;
  o_Energy_Bin_Pos_613  <= s_Energy_Bin_Pos_613  ;
  o_Energy_Bin_Pos_614  <= s_Energy_Bin_Pos_614  ;
  o_Energy_Bin_Pos_615  <= s_Energy_Bin_Pos_615  ;
  o_Energy_Bin_Pos_616  <= s_Energy_Bin_Pos_616  ;
  o_Energy_Bin_Pos_617  <= s_Energy_Bin_Pos_617  ;
  o_Energy_Bin_Pos_618  <= s_Energy_Bin_Pos_618  ;
  o_Energy_Bin_Pos_619  <= s_Energy_Bin_Pos_619  ;
  o_Energy_Bin_Pos_620  <= s_Energy_Bin_Pos_620  ;
  o_Energy_Bin_Pos_621  <= s_Energy_Bin_Pos_621  ;
  o_Energy_Bin_Pos_622  <= s_Energy_Bin_Pos_622  ;
  o_Energy_Bin_Pos_623  <= s_Energy_Bin_Pos_623  ;
  o_Energy_Bin_Pos_624  <= s_Energy_Bin_Pos_624  ;
  o_Energy_Bin_Pos_625  <= s_Energy_Bin_Pos_625  ;
  o_Energy_Bin_Pos_626  <= s_Energy_Bin_Pos_626  ;
  o_Energy_Bin_Pos_627  <= s_Energy_Bin_Pos_627  ;
  o_Energy_Bin_Pos_628  <= s_Energy_Bin_Pos_628  ;
  o_Energy_Bin_Pos_629  <= s_Energy_Bin_Pos_629  ;
  o_Energy_Bin_Pos_630  <= s_Energy_Bin_Pos_630  ;
  o_Energy_Bin_Pos_631  <= s_Energy_Bin_Pos_631  ;
  o_Energy_Bin_Pos_632  <= s_Energy_Bin_Pos_632  ;
  o_Energy_Bin_Pos_633  <= s_Energy_Bin_Pos_633  ;
  o_Energy_Bin_Pos_634  <= s_Energy_Bin_Pos_634  ;
  o_Energy_Bin_Pos_635  <= s_Energy_Bin_Pos_635  ;
  o_Energy_Bin_Pos_636  <= s_Energy_Bin_Pos_636  ;
  o_Energy_Bin_Pos_637  <= s_Energy_Bin_Pos_637  ;
  o_Energy_Bin_Pos_638  <= s_Energy_Bin_Pos_638  ;
  o_Energy_Bin_Pos_639  <= s_Energy_Bin_Pos_639  ;
  o_Energy_Bin_Pos_640  <= s_Energy_Bin_Pos_640  ;
  o_Energy_Bin_Pos_641  <= s_Energy_Bin_Pos_641  ;
  o_Energy_Bin_Pos_642  <= s_Energy_Bin_Pos_642  ;
  o_Energy_Bin_Pos_643  <= s_Energy_Bin_Pos_643  ;
  o_Energy_Bin_Pos_644  <= s_Energy_Bin_Pos_644  ;
  o_Energy_Bin_Pos_645  <= s_Energy_Bin_Pos_645  ;
  o_Energy_Bin_Pos_646  <= s_Energy_Bin_Pos_646  ;
  o_Energy_Bin_Pos_647  <= s_Energy_Bin_Pos_647  ;
  o_Energy_Bin_Pos_648  <= s_Energy_Bin_Pos_648  ;
  o_Energy_Bin_Pos_649  <= s_Energy_Bin_Pos_649  ;
  o_Energy_Bin_Pos_650  <= s_Energy_Bin_Pos_650  ;
  o_Energy_Bin_Pos_651  <= s_Energy_Bin_Pos_651  ;
  o_Energy_Bin_Pos_652  <= s_Energy_Bin_Pos_652  ;
  o_Energy_Bin_Pos_653  <= s_Energy_Bin_Pos_653  ;
  o_Energy_Bin_Pos_654  <= s_Energy_Bin_Pos_654  ;
  o_Energy_Bin_Pos_655  <= s_Energy_Bin_Pos_655  ;
  o_Energy_Bin_Pos_656  <= s_Energy_Bin_Pos_656  ;
  o_Energy_Bin_Pos_657  <= s_Energy_Bin_Pos_657  ;
  o_Energy_Bin_Pos_658  <= s_Energy_Bin_Pos_658  ;
  o_Energy_Bin_Pos_659  <= s_Energy_Bin_Pos_659  ;
  o_Energy_Bin_Pos_660  <= s_Energy_Bin_Pos_660  ;
  o_Energy_Bin_Pos_661  <= s_Energy_Bin_Pos_661  ;
  o_Energy_Bin_Pos_662  <= s_Energy_Bin_Pos_662  ;
  o_Energy_Bin_Pos_663  <= s_Energy_Bin_Pos_663  ;
  o_Energy_Bin_Pos_664  <= s_Energy_Bin_Pos_664  ;
  o_Energy_Bin_Pos_665  <= s_Energy_Bin_Pos_665  ;
  o_Energy_Bin_Pos_666  <= s_Energy_Bin_Pos_666  ;
  o_Energy_Bin_Pos_667  <= s_Energy_Bin_Pos_667  ;
  o_Energy_Bin_Pos_668  <= s_Energy_Bin_Pos_668  ;
  o_Energy_Bin_Pos_669  <= s_Energy_Bin_Pos_669  ;
  o_Energy_Bin_Pos_670  <= s_Energy_Bin_Pos_670  ;
  o_Energy_Bin_Pos_671  <= s_Energy_Bin_Pos_671  ;
  o_Energy_Bin_Pos_672  <= s_Energy_Bin_Pos_672  ;
  o_Energy_Bin_Pos_673  <= s_Energy_Bin_Pos_673  ;
  o_Energy_Bin_Pos_674  <= s_Energy_Bin_Pos_674  ;
  o_Energy_Bin_Pos_675  <= s_Energy_Bin_Pos_675  ;
  o_Energy_Bin_Pos_676  <= s_Energy_Bin_Pos_676  ;
  o_Energy_Bin_Pos_677  <= s_Energy_Bin_Pos_677  ;
  o_Energy_Bin_Pos_678  <= s_Energy_Bin_Pos_678  ;
  o_Energy_Bin_Pos_679  <= s_Energy_Bin_Pos_679  ;
  o_Energy_Bin_Pos_680  <= s_Energy_Bin_Pos_680  ;
  o_Energy_Bin_Pos_681  <= s_Energy_Bin_Pos_681  ;
  o_Energy_Bin_Pos_682  <= s_Energy_Bin_Pos_682  ;
  o_Energy_Bin_Pos_683  <= s_Energy_Bin_Pos_683  ;
  o_Energy_Bin_Pos_684  <= s_Energy_Bin_Pos_684  ;
  o_Energy_Bin_Pos_685  <= s_Energy_Bin_Pos_685  ;
  o_Energy_Bin_Pos_686  <= s_Energy_Bin_Pos_686  ;
  o_Energy_Bin_Pos_687  <= s_Energy_Bin_Pos_687  ;
  o_Energy_Bin_Pos_688  <= s_Energy_Bin_Pos_688  ;
  o_Energy_Bin_Pos_689  <= s_Energy_Bin_Pos_689  ;
  o_Energy_Bin_Pos_690  <= s_Energy_Bin_Pos_690  ;
  o_Energy_Bin_Pos_691  <= s_Energy_Bin_Pos_691  ;
  o_Energy_Bin_Pos_692  <= s_Energy_Bin_Pos_692  ;
  o_Energy_Bin_Pos_693  <= s_Energy_Bin_Pos_693  ;
  o_Energy_Bin_Pos_694  <= s_Energy_Bin_Pos_694  ;
  o_Energy_Bin_Pos_695  <= s_Energy_Bin_Pos_695  ;
  o_Energy_Bin_Pos_696  <= s_Energy_Bin_Pos_696  ;
  o_Energy_Bin_Pos_697  <= s_Energy_Bin_Pos_697  ;
  o_Energy_Bin_Pos_698  <= s_Energy_Bin_Pos_698  ;
  o_Energy_Bin_Pos_699  <= s_Energy_Bin_Pos_699  ;
  o_Energy_Bin_Pos_700  <= s_Energy_Bin_Pos_700  ;
  o_Energy_Bin_Pos_701  <= s_Energy_Bin_Pos_701  ;
  o_Energy_Bin_Pos_702  <= s_Energy_Bin_Pos_702  ;
  o_Energy_Bin_Pos_703  <= s_Energy_Bin_Pos_703  ;
  o_Energy_Bin_Pos_704  <= s_Energy_Bin_Pos_704  ;
  o_Energy_Bin_Pos_705  <= s_Energy_Bin_Pos_705  ;
  o_Energy_Bin_Pos_706  <= s_Energy_Bin_Pos_706  ;
  o_Energy_Bin_Pos_707  <= s_Energy_Bin_Pos_707  ;
  o_Energy_Bin_Pos_708  <= s_Energy_Bin_Pos_708  ;
  o_Energy_Bin_Pos_709  <= s_Energy_Bin_Pos_709  ;
  o_Energy_Bin_Pos_710  <= s_Energy_Bin_Pos_710  ;
  o_Energy_Bin_Pos_711  <= s_Energy_Bin_Pos_711  ;
  o_Energy_Bin_Pos_712  <= s_Energy_Bin_Pos_712  ;
  o_Energy_Bin_Pos_713  <= s_Energy_Bin_Pos_713  ;
  o_Energy_Bin_Pos_714  <= s_Energy_Bin_Pos_714  ;
  o_Energy_Bin_Pos_715  <= s_Energy_Bin_Pos_715  ;
  o_Energy_Bin_Pos_716  <= s_Energy_Bin_Pos_716  ;
  o_Energy_Bin_Pos_717  <= s_Energy_Bin_Pos_717  ;
  o_Energy_Bin_Pos_718  <= s_Energy_Bin_Pos_718  ;
  o_Energy_Bin_Pos_719  <= s_Energy_Bin_Pos_719  ;
  o_Energy_Bin_Pos_720  <= s_Energy_Bin_Pos_720  ;
  o_Energy_Bin_Pos_721  <= s_Energy_Bin_Pos_721  ;
  o_Energy_Bin_Pos_722  <= s_Energy_Bin_Pos_722  ;
  o_Energy_Bin_Pos_723  <= s_Energy_Bin_Pos_723  ;
  o_Energy_Bin_Pos_724  <= s_Energy_Bin_Pos_724  ;
  o_Energy_Bin_Pos_725  <= s_Energy_Bin_Pos_725  ;
  o_Energy_Bin_Pos_726  <= s_Energy_Bin_Pos_726  ;
  o_Energy_Bin_Pos_727  <= s_Energy_Bin_Pos_727  ;
  o_Energy_Bin_Pos_728  <= s_Energy_Bin_Pos_728  ;
  o_Energy_Bin_Pos_729  <= s_Energy_Bin_Pos_729  ;
  o_Energy_Bin_Pos_730  <= s_Energy_Bin_Pos_730  ;
  o_Energy_Bin_Pos_731  <= s_Energy_Bin_Pos_731  ;
  o_Energy_Bin_Pos_732  <= s_Energy_Bin_Pos_732  ;
  o_Energy_Bin_Pos_733  <= s_Energy_Bin_Pos_733  ;
  o_Energy_Bin_Pos_734  <= s_Energy_Bin_Pos_734  ;
  o_Energy_Bin_Pos_735  <= s_Energy_Bin_Pos_735  ;
  o_Energy_Bin_Pos_736  <= s_Energy_Bin_Pos_736  ;
  o_Energy_Bin_Pos_737  <= s_Energy_Bin_Pos_737  ;
  o_Energy_Bin_Pos_738  <= s_Energy_Bin_Pos_738  ;
  o_Energy_Bin_Pos_739  <= s_Energy_Bin_Pos_739  ;
  o_Energy_Bin_Pos_740  <= s_Energy_Bin_Pos_740  ;
  o_Energy_Bin_Pos_741  <= s_Energy_Bin_Pos_741  ;
  o_Energy_Bin_Pos_742  <= s_Energy_Bin_Pos_742  ;
  o_Energy_Bin_Pos_743  <= s_Energy_Bin_Pos_743  ;
  o_Energy_Bin_Pos_744  <= s_Energy_Bin_Pos_744  ;
  o_Energy_Bin_Pos_745  <= s_Energy_Bin_Pos_745  ;
  o_Energy_Bin_Pos_746  <= s_Energy_Bin_Pos_746  ;
  o_Energy_Bin_Pos_747  <= s_Energy_Bin_Pos_747  ;
  o_Energy_Bin_Pos_748  <= s_Energy_Bin_Pos_748  ;
  o_Energy_Bin_Pos_749  <= s_Energy_Bin_Pos_749  ;
  o_Energy_Bin_Pos_750  <= s_Energy_Bin_Pos_750  ;
  o_Energy_Bin_Pos_751  <= s_Energy_Bin_Pos_751  ;
  o_Energy_Bin_Pos_752  <= s_Energy_Bin_Pos_752  ;
  o_Energy_Bin_Pos_753  <= s_Energy_Bin_Pos_753  ;
  o_Energy_Bin_Pos_754  <= s_Energy_Bin_Pos_754  ;
  o_Energy_Bin_Pos_755  <= s_Energy_Bin_Pos_755  ;
  o_Energy_Bin_Pos_756  <= s_Energy_Bin_Pos_756  ;
  o_Energy_Bin_Pos_757  <= s_Energy_Bin_Pos_757  ;
  o_Energy_Bin_Pos_758  <= s_Energy_Bin_Pos_758  ;
  o_Energy_Bin_Pos_759  <= s_Energy_Bin_Pos_759  ;
  o_Energy_Bin_Pos_760  <= s_Energy_Bin_Pos_760  ;
  o_Energy_Bin_Pos_761  <= s_Energy_Bin_Pos_761  ;
  o_Energy_Bin_Pos_762  <= s_Energy_Bin_Pos_762  ;
  o_Energy_Bin_Pos_763  <= s_Energy_Bin_Pos_763  ;
  o_Energy_Bin_Pos_764  <= s_Energy_Bin_Pos_764  ;
  o_Energy_Bin_Pos_765  <= s_Energy_Bin_Pos_765  ;
  o_Energy_Bin_Pos_766  <= s_Energy_Bin_Pos_766  ;
  o_Energy_Bin_Pos_767  <= s_Energy_Bin_Pos_767  ;
  o_Energy_Bin_Pos_768  <= s_Energy_Bin_Pos_768  ;
  o_Energy_Bin_Pos_769  <= s_Energy_Bin_Pos_769  ;
  o_Energy_Bin_Pos_770  <= s_Energy_Bin_Pos_770  ;
  o_Energy_Bin_Pos_771  <= s_Energy_Bin_Pos_771  ;
  o_Energy_Bin_Pos_772  <= s_Energy_Bin_Pos_772  ;
  o_Energy_Bin_Pos_773  <= s_Energy_Bin_Pos_773  ;
  o_Energy_Bin_Pos_774  <= s_Energy_Bin_Pos_774  ;
  o_Energy_Bin_Pos_775  <= s_Energy_Bin_Pos_775  ;
  o_Energy_Bin_Pos_776  <= s_Energy_Bin_Pos_776  ;
  o_Energy_Bin_Pos_777  <= s_Energy_Bin_Pos_777  ;
  o_Energy_Bin_Pos_778  <= s_Energy_Bin_Pos_778  ;
  o_Energy_Bin_Pos_779  <= s_Energy_Bin_Pos_779  ;
  o_Energy_Bin_Pos_780  <= s_Energy_Bin_Pos_780  ;
  o_Energy_Bin_Pos_781  <= s_Energy_Bin_Pos_781  ;
  o_Energy_Bin_Pos_782  <= s_Energy_Bin_Pos_782  ;
  o_Energy_Bin_Pos_783  <= s_Energy_Bin_Pos_783  ;
  o_Energy_Bin_Pos_784  <= s_Energy_Bin_Pos_784  ;
  o_Energy_Bin_Pos_785  <= s_Energy_Bin_Pos_785  ;
  o_Energy_Bin_Pos_786  <= s_Energy_Bin_Pos_786  ;
  o_Energy_Bin_Pos_787  <= s_Energy_Bin_Pos_787  ;
  o_Energy_Bin_Pos_788  <= s_Energy_Bin_Pos_788  ;
  o_Energy_Bin_Pos_789  <= s_Energy_Bin_Pos_789  ;
  o_Energy_Bin_Pos_790  <= s_Energy_Bin_Pos_790  ;
  o_Energy_Bin_Pos_791  <= s_Energy_Bin_Pos_791  ;
  o_Energy_Bin_Pos_792  <= s_Energy_Bin_Pos_792  ;
  o_Energy_Bin_Pos_793  <= s_Energy_Bin_Pos_793  ;
  o_Energy_Bin_Pos_794  <= s_Energy_Bin_Pos_794  ;
  o_Energy_Bin_Pos_795  <= s_Energy_Bin_Pos_795  ;
  o_Energy_Bin_Pos_796  <= s_Energy_Bin_Pos_796  ;
  o_Energy_Bin_Pos_797  <= s_Energy_Bin_Pos_797  ;
  o_Energy_Bin_Pos_798  <= s_Energy_Bin_Pos_798  ;
  o_Energy_Bin_Pos_799  <= s_Energy_Bin_Pos_799  ;
  o_Energy_Bin_Pos_800  <= s_Energy_Bin_Pos_800  ;
  o_Energy_Bin_Pos_801  <= s_Energy_Bin_Pos_801  ;
  o_Energy_Bin_Pos_802  <= s_Energy_Bin_Pos_802  ;
  o_Energy_Bin_Pos_803  <= s_Energy_Bin_Pos_803  ;
  o_Energy_Bin_Pos_804  <= s_Energy_Bin_Pos_804  ;
  o_Energy_Bin_Pos_805  <= s_Energy_Bin_Pos_805  ;
  o_Energy_Bin_Pos_806  <= s_Energy_Bin_Pos_806  ;
  o_Energy_Bin_Pos_807  <= s_Energy_Bin_Pos_807  ;
  o_Energy_Bin_Pos_808  <= s_Energy_Bin_Pos_808  ;
  o_Energy_Bin_Pos_809  <= s_Energy_Bin_Pos_809  ;
  o_Energy_Bin_Pos_810  <= s_Energy_Bin_Pos_810  ;
  o_Energy_Bin_Pos_811  <= s_Energy_Bin_Pos_811  ;
  o_Energy_Bin_Pos_812  <= s_Energy_Bin_Pos_812  ;
  o_Energy_Bin_Pos_813  <= s_Energy_Bin_Pos_813  ;
  o_Energy_Bin_Pos_814  <= s_Energy_Bin_Pos_814  ;
  o_Energy_Bin_Pos_815  <= s_Energy_Bin_Pos_815  ;
  o_Energy_Bin_Pos_816  <= s_Energy_Bin_Pos_816  ;
  o_Energy_Bin_Pos_817  <= s_Energy_Bin_Pos_817  ;
  o_Energy_Bin_Pos_818  <= s_Energy_Bin_Pos_818  ;
  o_Energy_Bin_Pos_819  <= s_Energy_Bin_Pos_819  ;
  o_Energy_Bin_Pos_820  <= s_Energy_Bin_Pos_820  ;
  o_Energy_Bin_Pos_821  <= s_Energy_Bin_Pos_821  ;
  o_Energy_Bin_Pos_822  <= s_Energy_Bin_Pos_822  ;
  o_Energy_Bin_Pos_823  <= s_Energy_Bin_Pos_823  ;
  o_Energy_Bin_Pos_824  <= s_Energy_Bin_Pos_824  ;
  o_Energy_Bin_Pos_825  <= s_Energy_Bin_Pos_825  ;
  o_Energy_Bin_Pos_826  <= s_Energy_Bin_Pos_826  ;
  o_Energy_Bin_Pos_827  <= s_Energy_Bin_Pos_827  ;
  o_Energy_Bin_Pos_828  <= s_Energy_Bin_Pos_828  ;
  o_Energy_Bin_Pos_829  <= s_Energy_Bin_Pos_829  ;
  o_Energy_Bin_Pos_830  <= s_Energy_Bin_Pos_830  ;
  o_Energy_Bin_Pos_831  <= s_Energy_Bin_Pos_831  ;
  o_Energy_Bin_Pos_832  <= s_Energy_Bin_Pos_832  ;
  o_Energy_Bin_Pos_833  <= s_Energy_Bin_Pos_833  ;
  o_Energy_Bin_Pos_834  <= s_Energy_Bin_Pos_834  ;
  o_Energy_Bin_Pos_835  <= s_Energy_Bin_Pos_835  ;
  o_Energy_Bin_Pos_836  <= s_Energy_Bin_Pos_836  ;
  o_Energy_Bin_Pos_837  <= s_Energy_Bin_Pos_837  ;
  o_Energy_Bin_Pos_838  <= s_Energy_Bin_Pos_838  ;
  o_Energy_Bin_Pos_839  <= s_Energy_Bin_Pos_839  ;
  o_Energy_Bin_Pos_840  <= s_Energy_Bin_Pos_840  ;
  o_Energy_Bin_Pos_841  <= s_Energy_Bin_Pos_841  ;
  o_Energy_Bin_Pos_842  <= s_Energy_Bin_Pos_842  ;
  o_Energy_Bin_Pos_843  <= s_Energy_Bin_Pos_843  ;
  o_Energy_Bin_Pos_844  <= s_Energy_Bin_Pos_844  ;
  o_Energy_Bin_Pos_845  <= s_Energy_Bin_Pos_845  ;
  o_Energy_Bin_Pos_846  <= s_Energy_Bin_Pos_846  ;
  o_Energy_Bin_Pos_847  <= s_Energy_Bin_Pos_847  ;
  o_Energy_Bin_Pos_848  <= s_Energy_Bin_Pos_848  ;
  o_Energy_Bin_Pos_849  <= s_Energy_Bin_Pos_849  ;
  o_Energy_Bin_Pos_850  <= s_Energy_Bin_Pos_850  ;
  o_Energy_Bin_Pos_851  <= s_Energy_Bin_Pos_851  ;
  o_Energy_Bin_Pos_852  <= s_Energy_Bin_Pos_852  ;
  o_Energy_Bin_Pos_853  <= s_Energy_Bin_Pos_853  ;
  o_Energy_Bin_Pos_854  <= s_Energy_Bin_Pos_854  ;
  o_Energy_Bin_Pos_855  <= s_Energy_Bin_Pos_855  ;
  o_Energy_Bin_Pos_856  <= s_Energy_Bin_Pos_856  ;
  o_Energy_Bin_Pos_857  <= s_Energy_Bin_Pos_857  ;
  o_Energy_Bin_Pos_858  <= s_Energy_Bin_Pos_858  ;
  o_Energy_Bin_Pos_859  <= s_Energy_Bin_Pos_859  ;
  o_Energy_Bin_Pos_860  <= s_Energy_Bin_Pos_860  ;
  o_Energy_Bin_Pos_861  <= s_Energy_Bin_Pos_861  ;
  o_Energy_Bin_Pos_862  <= s_Energy_Bin_Pos_862  ;
  o_Energy_Bin_Pos_863  <= s_Energy_Bin_Pos_863  ;
  o_Energy_Bin_Pos_864  <= s_Energy_Bin_Pos_864  ;
  o_Energy_Bin_Pos_865  <= s_Energy_Bin_Pos_865  ;
  o_Energy_Bin_Pos_866  <= s_Energy_Bin_Pos_866  ;
  o_Energy_Bin_Pos_867  <= s_Energy_Bin_Pos_867  ;
  o_Energy_Bin_Pos_868  <= s_Energy_Bin_Pos_868  ;
  o_Energy_Bin_Pos_869  <= s_Energy_Bin_Pos_869  ;
  o_Energy_Bin_Pos_870  <= s_Energy_Bin_Pos_870  ;
  o_Energy_Bin_Pos_871  <= s_Energy_Bin_Pos_871  ;
  o_Energy_Bin_Pos_872  <= s_Energy_Bin_Pos_872  ;
  o_Energy_Bin_Pos_873  <= s_Energy_Bin_Pos_873  ;
  o_Energy_Bin_Pos_874  <= s_Energy_Bin_Pos_874  ;
  o_Energy_Bin_Pos_875  <= s_Energy_Bin_Pos_875  ;
  o_Energy_Bin_Pos_876  <= s_Energy_Bin_Pos_876  ;
  o_Energy_Bin_Pos_877  <= s_Energy_Bin_Pos_877  ;
  o_Energy_Bin_Pos_878  <= s_Energy_Bin_Pos_878  ;
  o_Energy_Bin_Pos_879  <= s_Energy_Bin_Pos_879  ;
  o_Energy_Bin_Pos_880  <= s_Energy_Bin_Pos_880  ;
  o_Energy_Bin_Pos_881  <= s_Energy_Bin_Pos_881  ;
  o_Energy_Bin_Pos_882  <= s_Energy_Bin_Pos_882  ;
  o_Energy_Bin_Pos_883  <= s_Energy_Bin_Pos_883  ;
  o_Energy_Bin_Pos_884  <= s_Energy_Bin_Pos_884  ;
  o_Energy_Bin_Pos_885  <= s_Energy_Bin_Pos_885  ;
  o_Energy_Bin_Pos_886  <= s_Energy_Bin_Pos_886  ;
  o_Energy_Bin_Pos_887  <= s_Energy_Bin_Pos_887  ;
  o_Energy_Bin_Pos_888  <= s_Energy_Bin_Pos_888  ;
  o_Energy_Bin_Pos_889  <= s_Energy_Bin_Pos_889  ;
  o_Energy_Bin_Pos_890  <= s_Energy_Bin_Pos_890  ;
  o_Energy_Bin_Pos_891  <= s_Energy_Bin_Pos_891  ;
  o_Energy_Bin_Pos_892  <= s_Energy_Bin_Pos_892  ;
  o_Energy_Bin_Pos_893  <= s_Energy_Bin_Pos_893  ;
  o_Energy_Bin_Pos_894  <= s_Energy_Bin_Pos_894  ;
  o_Energy_Bin_Pos_895  <= s_Energy_Bin_Pos_895  ;
  o_Energy_Bin_Pos_896  <= s_Energy_Bin_Pos_896  ;
  o_Energy_Bin_Pos_897  <= s_Energy_Bin_Pos_897  ;
  o_Energy_Bin_Pos_898  <= s_Energy_Bin_Pos_898  ;
  o_Energy_Bin_Pos_899  <= s_Energy_Bin_Pos_899  ;
  o_Energy_Bin_Pos_900  <= s_Energy_Bin_Pos_900  ;
  o_Energy_Bin_Pos_901  <= s_Energy_Bin_Pos_901  ;
  o_Energy_Bin_Pos_902  <= s_Energy_Bin_Pos_902  ;
  o_Energy_Bin_Pos_903  <= s_Energy_Bin_Pos_903  ;
  o_Energy_Bin_Pos_904  <= s_Energy_Bin_Pos_904  ;
  o_Energy_Bin_Pos_905  <= s_Energy_Bin_Pos_905  ;
  o_Energy_Bin_Pos_906  <= s_Energy_Bin_Pos_906  ;
  o_Energy_Bin_Pos_907  <= s_Energy_Bin_Pos_907  ;
  o_Energy_Bin_Pos_908  <= s_Energy_Bin_Pos_908  ;
  o_Energy_Bin_Pos_909  <= s_Energy_Bin_Pos_909  ;
  o_Energy_Bin_Pos_910  <= s_Energy_Bin_Pos_910  ;
  o_Energy_Bin_Pos_911  <= s_Energy_Bin_Pos_911  ;
  o_Energy_Bin_Pos_912  <= s_Energy_Bin_Pos_912  ;
  o_Energy_Bin_Pos_913  <= s_Energy_Bin_Pos_913  ;
  o_Energy_Bin_Pos_914  <= s_Energy_Bin_Pos_914  ;
  o_Energy_Bin_Pos_915  <= s_Energy_Bin_Pos_915  ;
  o_Energy_Bin_Pos_916  <= s_Energy_Bin_Pos_916  ;
  o_Energy_Bin_Pos_917  <= s_Energy_Bin_Pos_917  ;
  o_Energy_Bin_Pos_918  <= s_Energy_Bin_Pos_918  ;
  o_Energy_Bin_Pos_919  <= s_Energy_Bin_Pos_919  ;
  o_Energy_Bin_Pos_920  <= s_Energy_Bin_Pos_920  ;
  o_Energy_Bin_Pos_921  <= s_Energy_Bin_Pos_921  ;
  o_Energy_Bin_Pos_922  <= s_Energy_Bin_Pos_922  ;
  o_Energy_Bin_Pos_923  <= s_Energy_Bin_Pos_923  ;
  o_Energy_Bin_Pos_924  <= s_Energy_Bin_Pos_924  ;
  o_Energy_Bin_Pos_925  <= s_Energy_Bin_Pos_925  ;
  o_Energy_Bin_Pos_926  <= s_Energy_Bin_Pos_926  ;
  o_Energy_Bin_Pos_927  <= s_Energy_Bin_Pos_927  ;
  o_Energy_Bin_Pos_928  <= s_Energy_Bin_Pos_928  ;
  o_Energy_Bin_Pos_929  <= s_Energy_Bin_Pos_929  ;
  o_Energy_Bin_Pos_930  <= s_Energy_Bin_Pos_930  ;
  o_Energy_Bin_Pos_931  <= s_Energy_Bin_Pos_931  ;
  o_Energy_Bin_Pos_932  <= s_Energy_Bin_Pos_932  ;
  o_Energy_Bin_Pos_933  <= s_Energy_Bin_Pos_933  ;
  o_Energy_Bin_Pos_934  <= s_Energy_Bin_Pos_934  ;
  o_Energy_Bin_Pos_935  <= s_Energy_Bin_Pos_935  ;
  o_Energy_Bin_Pos_936  <= s_Energy_Bin_Pos_936  ;
  o_Energy_Bin_Pos_937  <= s_Energy_Bin_Pos_937  ;
  o_Energy_Bin_Pos_938  <= s_Energy_Bin_Pos_938  ;
  o_Energy_Bin_Pos_939  <= s_Energy_Bin_Pos_939  ;
  o_Energy_Bin_Pos_940  <= s_Energy_Bin_Pos_940  ;
  o_Energy_Bin_Pos_941  <= s_Energy_Bin_Pos_941  ;
  o_Energy_Bin_Pos_942  <= s_Energy_Bin_Pos_942  ;
  o_Energy_Bin_Pos_943  <= s_Energy_Bin_Pos_943  ;
  o_Energy_Bin_Pos_944  <= s_Energy_Bin_Pos_944  ;
  o_Energy_Bin_Pos_945  <= s_Energy_Bin_Pos_945  ;
  o_Energy_Bin_Pos_946  <= s_Energy_Bin_Pos_946  ;
  o_Energy_Bin_Pos_947  <= s_Energy_Bin_Pos_947  ;
  o_Energy_Bin_Pos_948  <= s_Energy_Bin_Pos_948  ;
  o_Energy_Bin_Pos_949  <= s_Energy_Bin_Pos_949  ;
  o_Energy_Bin_Pos_950  <= s_Energy_Bin_Pos_950  ;
  o_Energy_Bin_Pos_951  <= s_Energy_Bin_Pos_951  ;
  o_Energy_Bin_Pos_952  <= s_Energy_Bin_Pos_952  ;
  o_Energy_Bin_Pos_953  <= s_Energy_Bin_Pos_953  ;
  o_Energy_Bin_Pos_954  <= s_Energy_Bin_Pos_954  ;
  o_Energy_Bin_Pos_955  <= s_Energy_Bin_Pos_955  ;
  o_Energy_Bin_Pos_956  <= s_Energy_Bin_Pos_956  ;
  o_Energy_Bin_Pos_957  <= s_Energy_Bin_Pos_957  ;
  o_Energy_Bin_Pos_958  <= s_Energy_Bin_Pos_958  ;
  o_Energy_Bin_Pos_959  <= s_Energy_Bin_Pos_959  ;
  o_Energy_Bin_Pos_960  <= s_Energy_Bin_Pos_960  ;
  o_Energy_Bin_Pos_961  <= s_Energy_Bin_Pos_961  ;
  o_Energy_Bin_Pos_962  <= s_Energy_Bin_Pos_962  ;
  o_Energy_Bin_Pos_963  <= s_Energy_Bin_Pos_963  ;
  o_Energy_Bin_Pos_964  <= s_Energy_Bin_Pos_964  ;
  o_Energy_Bin_Pos_965  <= s_Energy_Bin_Pos_965  ;
  o_Energy_Bin_Pos_966  <= s_Energy_Bin_Pos_966  ;
  o_Energy_Bin_Pos_967  <= s_Energy_Bin_Pos_967  ;
  o_Energy_Bin_Pos_968  <= s_Energy_Bin_Pos_968  ;
  o_Energy_Bin_Pos_969  <= s_Energy_Bin_Pos_969  ;
  o_Energy_Bin_Pos_970  <= s_Energy_Bin_Pos_970  ;
  o_Energy_Bin_Pos_971  <= s_Energy_Bin_Pos_971  ;
  o_Energy_Bin_Pos_972  <= s_Energy_Bin_Pos_972  ;
  o_Energy_Bin_Pos_973  <= s_Energy_Bin_Pos_973  ;
  o_Energy_Bin_Pos_974  <= s_Energy_Bin_Pos_974  ;
  o_Energy_Bin_Pos_975  <= s_Energy_Bin_Pos_975  ;
  o_Energy_Bin_Pos_976  <= s_Energy_Bin_Pos_976  ;
  o_Energy_Bin_Pos_977  <= s_Energy_Bin_Pos_977  ;
  o_Energy_Bin_Pos_978  <= s_Energy_Bin_Pos_978  ;
  o_Energy_Bin_Pos_979  <= s_Energy_Bin_Pos_979  ;
  o_Energy_Bin_Pos_980  <= s_Energy_Bin_Pos_980  ;
  o_Energy_Bin_Pos_981  <= s_Energy_Bin_Pos_981  ;
  o_Energy_Bin_Pos_982  <= s_Energy_Bin_Pos_982  ;
  o_Energy_Bin_Pos_983  <= s_Energy_Bin_Pos_983  ;
  o_Energy_Bin_Pos_984  <= s_Energy_Bin_Pos_984  ;
  o_Energy_Bin_Pos_985  <= s_Energy_Bin_Pos_985  ;
  o_Energy_Bin_Pos_986  <= s_Energy_Bin_Pos_986  ;
  o_Energy_Bin_Pos_987  <= s_Energy_Bin_Pos_987  ;
  o_Energy_Bin_Pos_988  <= s_Energy_Bin_Pos_988  ;
  o_Energy_Bin_Pos_989  <= s_Energy_Bin_Pos_989  ;
  o_Energy_Bin_Pos_990  <= s_Energy_Bin_Pos_990  ;
  o_Energy_Bin_Pos_991  <= s_Energy_Bin_Pos_991  ;
  o_Energy_Bin_Pos_992  <= s_Energy_Bin_Pos_992  ;
  o_Energy_Bin_Pos_993  <= s_Energy_Bin_Pos_993  ;
  o_Energy_Bin_Pos_994  <= s_Energy_Bin_Pos_994  ;
  o_Energy_Bin_Pos_995  <= s_Energy_Bin_Pos_995  ;
  o_Energy_Bin_Pos_996  <= s_Energy_Bin_Pos_996  ;
  o_Energy_Bin_Pos_997  <= s_Energy_Bin_Pos_997  ;
  o_Energy_Bin_Pos_998  <= s_Energy_Bin_Pos_998  ;
  o_Energy_Bin_Pos_999  <= s_Energy_Bin_Pos_999  ;
  o_Energy_Bin_Pos_1000 <= s_Energy_Bin_Pos_1000 ;
  o_Energy_Bin_Pos_1001 <= s_Energy_Bin_Pos_1001 ;
  o_Energy_Bin_Pos_1002 <= s_Energy_Bin_Pos_1002 ;
  o_Energy_Bin_Pos_1003 <= s_Energy_Bin_Pos_1003 ;
  o_Energy_Bin_Pos_1004 <= s_Energy_Bin_Pos_1004 ;
  o_Energy_Bin_Pos_1005 <= s_Energy_Bin_Pos_1005 ;
  o_Energy_Bin_Pos_1006 <= s_Energy_Bin_Pos_1006 ;
  o_Energy_Bin_Pos_1007 <= s_Energy_Bin_Pos_1007 ;
  o_Energy_Bin_Pos_1008 <= s_Energy_Bin_Pos_1008 ;
  o_Energy_Bin_Pos_1009 <= s_Energy_Bin_Pos_1009 ;
  o_Energy_Bin_Pos_1010 <= s_Energy_Bin_Pos_1010 ;
  o_Energy_Bin_Pos_1011 <= s_Energy_Bin_Pos_1011 ;
  o_Energy_Bin_Pos_1012 <= s_Energy_Bin_Pos_1012 ;
  o_Energy_Bin_Pos_1013 <= s_Energy_Bin_Pos_1013 ;
  o_Energy_Bin_Pos_1014 <= s_Energy_Bin_Pos_1014 ;
  o_Energy_Bin_Pos_1015 <= s_Energy_Bin_Pos_1015 ;
  o_Energy_Bin_Pos_1016 <= s_Energy_Bin_Pos_1016 ;
  o_Energy_Bin_Pos_1017 <= s_Energy_Bin_Pos_1017 ;
  o_Energy_Bin_Pos_1018 <= s_Energy_Bin_Pos_1018 ;
  o_Energy_Bin_Pos_1019 <= s_Energy_Bin_Pos_1019 ;
  o_Energy_Bin_Pos_1020 <= s_Energy_Bin_Pos_1020 ;
  o_Energy_Bin_Pos_1021 <= s_Energy_Bin_Pos_1021 ;
  o_Energy_Bin_Pos_1022 <= s_Energy_Bin_Pos_1022 ;
  o_Energy_Bin_Pos_1023 <= s_Energy_Bin_Pos_1023 ;
  o_Energy_Bin_Pos_1024 <= s_Energy_Bin_Pos_1024 ;
  
  
  o_Energy_Bin_1    <= s_Energy_Bin_1    ;
  o_Energy_Bin_2    <= s_Energy_Bin_2    ;
  o_Energy_Bin_3    <= s_Energy_Bin_3    ;
  o_Energy_Bin_4    <= s_Energy_Bin_4    ;
  o_Energy_Bin_5    <= s_Energy_Bin_5    ;
  o_Energy_Bin_6    <= s_Energy_Bin_6    ;
  o_Energy_Bin_7    <= s_Energy_Bin_7    ;
  o_Energy_Bin_8    <= s_Energy_Bin_8    ;
  o_Energy_Bin_9    <= s_Energy_Bin_9    ;
  o_Energy_Bin_10   <= s_Energy_Bin_10   ;
  o_Energy_Bin_11   <= s_Energy_Bin_11   ;
  o_Energy_Bin_12   <= s_Energy_Bin_12   ;
  o_Energy_Bin_13   <= s_Energy_Bin_13   ;
  o_Energy_Bin_14   <= s_Energy_Bin_14   ;
  o_Energy_Bin_15   <= s_Energy_Bin_15   ;
  o_Energy_Bin_16   <= s_Energy_Bin_16   ;
  o_Energy_Bin_17   <= s_Energy_Bin_17   ;
  o_Energy_Bin_18   <= s_Energy_Bin_18   ;
  o_Energy_Bin_19   <= s_Energy_Bin_19   ;
  o_Energy_Bin_20   <= s_Energy_Bin_20   ;
  o_Energy_Bin_21   <= s_Energy_Bin_21   ;
  o_Energy_Bin_22   <= s_Energy_Bin_22   ;
  o_Energy_Bin_23   <= s_Energy_Bin_23   ;
  o_Energy_Bin_24   <= s_Energy_Bin_24   ;
  o_Energy_Bin_25   <= s_Energy_Bin_25   ;
  o_Energy_Bin_26   <= s_Energy_Bin_26   ;
  o_Energy_Bin_27   <= s_Energy_Bin_27   ;
  o_Energy_Bin_28   <= s_Energy_Bin_28   ;
  o_Energy_Bin_29   <= s_Energy_Bin_29   ;
  o_Energy_Bin_30   <= s_Energy_Bin_30   ;
  o_Energy_Bin_31   <= s_Energy_Bin_31   ;
  o_Energy_Bin_32   <= s_Energy_Bin_32   ;
  o_Energy_Bin_33   <= s_Energy_Bin_33   ;
  o_Energy_Bin_34   <= s_Energy_Bin_34   ;
  o_Energy_Bin_35   <= s_Energy_Bin_35   ;
  o_Energy_Bin_36   <= s_Energy_Bin_36   ;
  o_Energy_Bin_37   <= s_Energy_Bin_37   ;
  o_Energy_Bin_38   <= s_Energy_Bin_38   ;
  o_Energy_Bin_39   <= s_Energy_Bin_39   ;
  o_Energy_Bin_40   <= s_Energy_Bin_40   ;
  o_Energy_Bin_41   <= s_Energy_Bin_41   ;
  o_Energy_Bin_42   <= s_Energy_Bin_42   ;
  o_Energy_Bin_43   <= s_Energy_Bin_43   ;
  o_Energy_Bin_44   <= s_Energy_Bin_44   ;
  o_Energy_Bin_45   <= s_Energy_Bin_45   ;
  o_Energy_Bin_46   <= s_Energy_Bin_46   ;
  o_Energy_Bin_47   <= s_Energy_Bin_47   ;
  o_Energy_Bin_48   <= s_Energy_Bin_48   ;
  o_Energy_Bin_49   <= s_Energy_Bin_49   ;
  o_Energy_Bin_50   <= s_Energy_Bin_50   ;
  o_Energy_Bin_51   <= s_Energy_Bin_51   ;
  o_Energy_Bin_52   <= s_Energy_Bin_52   ;
  o_Energy_Bin_53   <= s_Energy_Bin_53   ;
  o_Energy_Bin_54   <= s_Energy_Bin_54   ;
  o_Energy_Bin_55   <= s_Energy_Bin_55   ;
  o_Energy_Bin_56   <= s_Energy_Bin_56   ;
  o_Energy_Bin_57   <= s_Energy_Bin_57   ;
  o_Energy_Bin_58   <= s_Energy_Bin_58   ;
  o_Energy_Bin_59   <= s_Energy_Bin_59   ;
  o_Energy_Bin_60   <= s_Energy_Bin_60   ;
  o_Energy_Bin_61   <= s_Energy_Bin_61   ;
  o_Energy_Bin_62   <= s_Energy_Bin_62   ;
  o_Energy_Bin_63   <= s_Energy_Bin_63   ;
  o_Energy_Bin_64   <= s_Energy_Bin_64   ;
  o_Energy_Bin_65   <= s_Energy_Bin_65   ;
  o_Energy_Bin_66   <= s_Energy_Bin_66   ;
  o_Energy_Bin_67   <= s_Energy_Bin_67   ;
  o_Energy_Bin_68   <= s_Energy_Bin_68   ;
  o_Energy_Bin_69   <= s_Energy_Bin_69   ;
  o_Energy_Bin_70   <= s_Energy_Bin_70   ;
  o_Energy_Bin_71   <= s_Energy_Bin_71   ;
  o_Energy_Bin_72   <= s_Energy_Bin_72   ;
  o_Energy_Bin_73   <= s_Energy_Bin_73   ;
  o_Energy_Bin_74   <= s_Energy_Bin_74   ;
  o_Energy_Bin_75   <= s_Energy_Bin_75   ;
  o_Energy_Bin_76   <= s_Energy_Bin_76   ;
  o_Energy_Bin_77   <= s_Energy_Bin_77   ;
  o_Energy_Bin_78   <= s_Energy_Bin_78   ;
  o_Energy_Bin_79   <= s_Energy_Bin_79   ;
  o_Energy_Bin_80   <= s_Energy_Bin_80   ;
  o_Energy_Bin_81   <= s_Energy_Bin_81   ;
  o_Energy_Bin_82   <= s_Energy_Bin_82   ;
  o_Energy_Bin_83   <= s_Energy_Bin_83   ;
  o_Energy_Bin_84   <= s_Energy_Bin_84   ;
  o_Energy_Bin_85   <= s_Energy_Bin_85   ;
  o_Energy_Bin_86   <= s_Energy_Bin_86   ;
  o_Energy_Bin_87   <= s_Energy_Bin_87   ;
  o_Energy_Bin_88   <= s_Energy_Bin_88   ;
  o_Energy_Bin_89   <= s_Energy_Bin_89   ;
  o_Energy_Bin_90   <= s_Energy_Bin_90   ;
  o_Energy_Bin_91   <= s_Energy_Bin_91   ;
  o_Energy_Bin_92   <= s_Energy_Bin_92   ;
  o_Energy_Bin_93   <= s_Energy_Bin_93   ;
  o_Energy_Bin_94   <= s_Energy_Bin_94   ;
  o_Energy_Bin_95   <= s_Energy_Bin_95   ;
  o_Energy_Bin_96   <= s_Energy_Bin_96   ;
  o_Energy_Bin_97   <= s_Energy_Bin_97   ;
  o_Energy_Bin_98   <= s_Energy_Bin_98   ;
  o_Energy_Bin_99   <= s_Energy_Bin_99   ;
  o_Energy_Bin_100  <= s_Energy_Bin_100  ;
  o_Energy_Bin_101  <= s_Energy_Bin_101  ;
  o_Energy_Bin_102  <= s_Energy_Bin_102  ;
  o_Energy_Bin_103  <= s_Energy_Bin_103  ;
  o_Energy_Bin_104  <= s_Energy_Bin_104  ;
  o_Energy_Bin_105  <= s_Energy_Bin_105  ;
  o_Energy_Bin_106  <= s_Energy_Bin_106  ;
  o_Energy_Bin_107  <= s_Energy_Bin_107  ;
  o_Energy_Bin_108  <= s_Energy_Bin_108  ;
  o_Energy_Bin_109  <= s_Energy_Bin_109  ;
  o_Energy_Bin_110  <= s_Energy_Bin_110  ;
  o_Energy_Bin_111  <= s_Energy_Bin_111  ;
  o_Energy_Bin_112  <= s_Energy_Bin_112  ;
  o_Energy_Bin_113  <= s_Energy_Bin_113  ;
  o_Energy_Bin_114  <= s_Energy_Bin_114  ;
  o_Energy_Bin_115  <= s_Energy_Bin_115  ;
  o_Energy_Bin_116  <= s_Energy_Bin_116  ;
  o_Energy_Bin_117  <= s_Energy_Bin_117  ;
  o_Energy_Bin_118  <= s_Energy_Bin_118  ;
  o_Energy_Bin_119  <= s_Energy_Bin_119  ;
  o_Energy_Bin_120  <= s_Energy_Bin_120  ;
  o_Energy_Bin_121  <= s_Energy_Bin_121  ;
  o_Energy_Bin_122  <= s_Energy_Bin_122  ;
  o_Energy_Bin_123  <= s_Energy_Bin_123  ;
  o_Energy_Bin_124  <= s_Energy_Bin_124  ;
  o_Energy_Bin_125  <= s_Energy_Bin_125  ;
  o_Energy_Bin_126  <= s_Energy_Bin_126  ;
  o_Energy_Bin_127  <= s_Energy_Bin_127  ;
  o_Energy_Bin_128  <= s_Energy_Bin_128  ;
  o_Energy_Bin_129  <= s_Energy_Bin_129  ;
  o_Energy_Bin_130  <= s_Energy_Bin_130  ;
  o_Energy_Bin_131  <= s_Energy_Bin_131  ;
  o_Energy_Bin_132  <= s_Energy_Bin_132  ;
  o_Energy_Bin_133  <= s_Energy_Bin_133  ;
  o_Energy_Bin_134  <= s_Energy_Bin_134  ;
  o_Energy_Bin_135  <= s_Energy_Bin_135  ;
  o_Energy_Bin_136  <= s_Energy_Bin_136  ;
  o_Energy_Bin_137  <= s_Energy_Bin_137  ;
  o_Energy_Bin_138  <= s_Energy_Bin_138  ;
  o_Energy_Bin_139  <= s_Energy_Bin_139  ;
  o_Energy_Bin_140  <= s_Energy_Bin_140  ;
  o_Energy_Bin_141  <= s_Energy_Bin_141  ;
  o_Energy_Bin_142  <= s_Energy_Bin_142  ;
  o_Energy_Bin_143  <= s_Energy_Bin_143  ;
  o_Energy_Bin_144  <= s_Energy_Bin_144  ;
  o_Energy_Bin_145  <= s_Energy_Bin_145  ;
  o_Energy_Bin_146  <= s_Energy_Bin_146  ;
  o_Energy_Bin_147  <= s_Energy_Bin_147  ;
  o_Energy_Bin_148  <= s_Energy_Bin_148  ;
  o_Energy_Bin_149  <= s_Energy_Bin_149  ;
  o_Energy_Bin_150  <= s_Energy_Bin_150  ;
  o_Energy_Bin_151  <= s_Energy_Bin_151  ;
  o_Energy_Bin_152  <= s_Energy_Bin_152  ;
  o_Energy_Bin_153  <= s_Energy_Bin_153  ;
  o_Energy_Bin_154  <= s_Energy_Bin_154  ;
  o_Energy_Bin_155  <= s_Energy_Bin_155  ;
  o_Energy_Bin_156  <= s_Energy_Bin_156  ;
  o_Energy_Bin_157  <= s_Energy_Bin_157  ;
  o_Energy_Bin_158  <= s_Energy_Bin_158  ;
  o_Energy_Bin_159  <= s_Energy_Bin_159  ;
  o_Energy_Bin_160  <= s_Energy_Bin_160  ;
  o_Energy_Bin_161  <= s_Energy_Bin_161  ;
  o_Energy_Bin_162  <= s_Energy_Bin_162  ;
  o_Energy_Bin_163  <= s_Energy_Bin_163  ;
  o_Energy_Bin_164  <= s_Energy_Bin_164  ;
  o_Energy_Bin_165  <= s_Energy_Bin_165  ;
  o_Energy_Bin_166  <= s_Energy_Bin_166  ;
  o_Energy_Bin_167  <= s_Energy_Bin_167  ;
  o_Energy_Bin_168  <= s_Energy_Bin_168  ;
  o_Energy_Bin_169  <= s_Energy_Bin_169  ;
  o_Energy_Bin_170  <= s_Energy_Bin_170  ;
  o_Energy_Bin_171  <= s_Energy_Bin_171  ;
  o_Energy_Bin_172  <= s_Energy_Bin_172  ;
  o_Energy_Bin_173  <= s_Energy_Bin_173  ;
  o_Energy_Bin_174  <= s_Energy_Bin_174  ;
  o_Energy_Bin_175  <= s_Energy_Bin_175  ;
  o_Energy_Bin_176  <= s_Energy_Bin_176  ;
  o_Energy_Bin_177  <= s_Energy_Bin_177  ;
  o_Energy_Bin_178  <= s_Energy_Bin_178  ;
  o_Energy_Bin_179  <= s_Energy_Bin_179  ;
  o_Energy_Bin_180  <= s_Energy_Bin_180  ;
  o_Energy_Bin_181  <= s_Energy_Bin_181  ;
  o_Energy_Bin_182  <= s_Energy_Bin_182  ;
  o_Energy_Bin_183  <= s_Energy_Bin_183  ;
  o_Energy_Bin_184  <= s_Energy_Bin_184  ;
  o_Energy_Bin_185  <= s_Energy_Bin_185  ;
  o_Energy_Bin_186  <= s_Energy_Bin_186  ;
  o_Energy_Bin_187  <= s_Energy_Bin_187  ;
  o_Energy_Bin_188  <= s_Energy_Bin_188  ;
  o_Energy_Bin_189  <= s_Energy_Bin_189  ;
  o_Energy_Bin_190  <= s_Energy_Bin_190  ;
  o_Energy_Bin_191  <= s_Energy_Bin_191  ;
  o_Energy_Bin_192  <= s_Energy_Bin_192  ;
  o_Energy_Bin_193  <= s_Energy_Bin_193  ;
  o_Energy_Bin_194  <= s_Energy_Bin_194  ;
  o_Energy_Bin_195  <= s_Energy_Bin_195  ;
  o_Energy_Bin_196  <= s_Energy_Bin_196  ;
  o_Energy_Bin_197  <= s_Energy_Bin_197  ;
  o_Energy_Bin_198  <= s_Energy_Bin_198  ;
  o_Energy_Bin_199  <= s_Energy_Bin_199  ;
  o_Energy_Bin_200  <= s_Energy_Bin_200  ;
  o_Energy_Bin_201  <= s_Energy_Bin_201  ;
  o_Energy_Bin_202  <= s_Energy_Bin_202  ;
  o_Energy_Bin_203  <= s_Energy_Bin_203  ;
  o_Energy_Bin_204  <= s_Energy_Bin_204  ;
  o_Energy_Bin_205  <= s_Energy_Bin_205  ;
  o_Energy_Bin_206  <= s_Energy_Bin_206  ;
  o_Energy_Bin_207  <= s_Energy_Bin_207  ;
  o_Energy_Bin_208  <= s_Energy_Bin_208  ;
  o_Energy_Bin_209  <= s_Energy_Bin_209  ;
  o_Energy_Bin_210  <= s_Energy_Bin_210  ;
  o_Energy_Bin_211  <= s_Energy_Bin_211  ;
  o_Energy_Bin_212  <= s_Energy_Bin_212  ;
  o_Energy_Bin_213  <= s_Energy_Bin_213  ;
  o_Energy_Bin_214  <= s_Energy_Bin_214  ;
  o_Energy_Bin_215  <= s_Energy_Bin_215  ;
  o_Energy_Bin_216  <= s_Energy_Bin_216  ;
  o_Energy_Bin_217  <= s_Energy_Bin_217  ;
  o_Energy_Bin_218  <= s_Energy_Bin_218  ;
  o_Energy_Bin_219  <= s_Energy_Bin_219  ;
  o_Energy_Bin_220  <= s_Energy_Bin_220  ;
  o_Energy_Bin_221  <= s_Energy_Bin_221  ;
  o_Energy_Bin_222  <= s_Energy_Bin_222  ;
  o_Energy_Bin_223  <= s_Energy_Bin_223  ;
  o_Energy_Bin_224  <= s_Energy_Bin_224  ;
  o_Energy_Bin_225  <= s_Energy_Bin_225  ;
  o_Energy_Bin_226  <= s_Energy_Bin_226  ;
  o_Energy_Bin_227  <= s_Energy_Bin_227  ;
  o_Energy_Bin_228  <= s_Energy_Bin_228  ;
  o_Energy_Bin_229  <= s_Energy_Bin_229  ;
  o_Energy_Bin_230  <= s_Energy_Bin_230  ;
  o_Energy_Bin_231  <= s_Energy_Bin_231  ;
  o_Energy_Bin_232  <= s_Energy_Bin_232  ;
  o_Energy_Bin_233  <= s_Energy_Bin_233  ;
  o_Energy_Bin_234  <= s_Energy_Bin_234  ;
  o_Energy_Bin_235  <= s_Energy_Bin_235  ;
  o_Energy_Bin_236  <= s_Energy_Bin_236  ;
  o_Energy_Bin_237  <= s_Energy_Bin_237  ;
  o_Energy_Bin_238  <= s_Energy_Bin_238  ;
  o_Energy_Bin_239  <= s_Energy_Bin_239  ;
  o_Energy_Bin_240  <= s_Energy_Bin_240  ;
  o_Energy_Bin_241  <= s_Energy_Bin_241  ;
  o_Energy_Bin_242  <= s_Energy_Bin_242  ;
  o_Energy_Bin_243  <= s_Energy_Bin_243  ;
  o_Energy_Bin_244  <= s_Energy_Bin_244  ;
  o_Energy_Bin_245  <= s_Energy_Bin_245  ;
  o_Energy_Bin_246  <= s_Energy_Bin_246  ;
  o_Energy_Bin_247  <= s_Energy_Bin_247  ;
  o_Energy_Bin_248  <= s_Energy_Bin_248  ;
  o_Energy_Bin_249  <= s_Energy_Bin_249  ;
  o_Energy_Bin_250  <= s_Energy_Bin_250  ;
  o_Energy_Bin_251  <= s_Energy_Bin_251  ;
  o_Energy_Bin_252  <= s_Energy_Bin_252  ;
  o_Energy_Bin_253  <= s_Energy_Bin_253  ;
  o_Energy_Bin_254  <= s_Energy_Bin_254  ;
  o_Energy_Bin_255  <= s_Energy_Bin_255  ;
  o_Energy_Bin_256  <= s_Energy_Bin_256  ;
  o_Energy_Bin_257  <= s_Energy_Bin_257  ;
  o_Energy_Bin_258  <= s_Energy_Bin_258  ;
  o_Energy_Bin_259  <= s_Energy_Bin_259  ;
  o_Energy_Bin_260  <= s_Energy_Bin_260  ;
  o_Energy_Bin_261  <= s_Energy_Bin_261  ;
  o_Energy_Bin_262  <= s_Energy_Bin_262  ;
  o_Energy_Bin_263  <= s_Energy_Bin_263  ;
  o_Energy_Bin_264  <= s_Energy_Bin_264  ;
  o_Energy_Bin_265  <= s_Energy_Bin_265  ;
  o_Energy_Bin_266  <= s_Energy_Bin_266  ;
  o_Energy_Bin_267  <= s_Energy_Bin_267  ;
  o_Energy_Bin_268  <= s_Energy_Bin_268  ;
  o_Energy_Bin_269  <= s_Energy_Bin_269  ;
  o_Energy_Bin_270  <= s_Energy_Bin_270  ;
  o_Energy_Bin_271  <= s_Energy_Bin_271  ;
  o_Energy_Bin_272  <= s_Energy_Bin_272  ;
  o_Energy_Bin_273  <= s_Energy_Bin_273  ;
  o_Energy_Bin_274  <= s_Energy_Bin_274  ;
  o_Energy_Bin_275  <= s_Energy_Bin_275  ;
  o_Energy_Bin_276  <= s_Energy_Bin_276  ;
  o_Energy_Bin_277  <= s_Energy_Bin_277  ;
  o_Energy_Bin_278  <= s_Energy_Bin_278  ;
  o_Energy_Bin_279  <= s_Energy_Bin_279  ;
  o_Energy_Bin_280  <= s_Energy_Bin_280  ;
  o_Energy_Bin_281  <= s_Energy_Bin_281  ;
  o_Energy_Bin_282  <= s_Energy_Bin_282  ;
  o_Energy_Bin_283  <= s_Energy_Bin_283  ;
  o_Energy_Bin_284  <= s_Energy_Bin_284  ;
  o_Energy_Bin_285  <= s_Energy_Bin_285  ;
  o_Energy_Bin_286  <= s_Energy_Bin_286  ;
  o_Energy_Bin_287  <= s_Energy_Bin_287  ;
  o_Energy_Bin_288  <= s_Energy_Bin_288  ;
  o_Energy_Bin_289  <= s_Energy_Bin_289  ;
  o_Energy_Bin_290  <= s_Energy_Bin_290  ;
  o_Energy_Bin_291  <= s_Energy_Bin_291  ;
  o_Energy_Bin_292  <= s_Energy_Bin_292  ;
  o_Energy_Bin_293  <= s_Energy_Bin_293  ;
  o_Energy_Bin_294  <= s_Energy_Bin_294  ;
  o_Energy_Bin_295  <= s_Energy_Bin_295  ;
  o_Energy_Bin_296  <= s_Energy_Bin_296  ;
  o_Energy_Bin_297  <= s_Energy_Bin_297  ;
  o_Energy_Bin_298  <= s_Energy_Bin_298  ;
  o_Energy_Bin_299  <= s_Energy_Bin_299  ;
  o_Energy_Bin_300  <= s_Energy_Bin_300  ;
  o_Energy_Bin_301  <= s_Energy_Bin_301  ;
  o_Energy_Bin_302  <= s_Energy_Bin_302  ;
  o_Energy_Bin_303  <= s_Energy_Bin_303  ;
  o_Energy_Bin_304  <= s_Energy_Bin_304  ;
  o_Energy_Bin_305  <= s_Energy_Bin_305  ;
  o_Energy_Bin_306  <= s_Energy_Bin_306  ;
  o_Energy_Bin_307  <= s_Energy_Bin_307  ;
  o_Energy_Bin_308  <= s_Energy_Bin_308  ;
  o_Energy_Bin_309  <= s_Energy_Bin_309  ;
  o_Energy_Bin_310  <= s_Energy_Bin_310  ;
  o_Energy_Bin_311  <= s_Energy_Bin_311  ;
  o_Energy_Bin_312  <= s_Energy_Bin_312  ;
  o_Energy_Bin_313  <= s_Energy_Bin_313  ;
  o_Energy_Bin_314  <= s_Energy_Bin_314  ;
  o_Energy_Bin_315  <= s_Energy_Bin_315  ;
  o_Energy_Bin_316  <= s_Energy_Bin_316  ;
  o_Energy_Bin_317  <= s_Energy_Bin_317  ;
  o_Energy_Bin_318  <= s_Energy_Bin_318  ;
  o_Energy_Bin_319  <= s_Energy_Bin_319  ;
  o_Energy_Bin_320  <= s_Energy_Bin_320  ;
  o_Energy_Bin_321  <= s_Energy_Bin_321  ;
  o_Energy_Bin_322  <= s_Energy_Bin_322  ;
  o_Energy_Bin_323  <= s_Energy_Bin_323  ;
  o_Energy_Bin_324  <= s_Energy_Bin_324  ;
  o_Energy_Bin_325  <= s_Energy_Bin_325  ;
  o_Energy_Bin_326  <= s_Energy_Bin_326  ;
  o_Energy_Bin_327  <= s_Energy_Bin_327  ;
  o_Energy_Bin_328  <= s_Energy_Bin_328  ;
  o_Energy_Bin_329  <= s_Energy_Bin_329  ;
  o_Energy_Bin_330  <= s_Energy_Bin_330  ;
  o_Energy_Bin_331  <= s_Energy_Bin_331  ;
  o_Energy_Bin_332  <= s_Energy_Bin_332  ;
  o_Energy_Bin_333  <= s_Energy_Bin_333  ;
  o_Energy_Bin_334  <= s_Energy_Bin_334  ;
  o_Energy_Bin_335  <= s_Energy_Bin_335  ;
  o_Energy_Bin_336  <= s_Energy_Bin_336  ;
  o_Energy_Bin_337  <= s_Energy_Bin_337  ;
  o_Energy_Bin_338  <= s_Energy_Bin_338  ;
  o_Energy_Bin_339  <= s_Energy_Bin_339  ;
  o_Energy_Bin_340  <= s_Energy_Bin_340  ;
  o_Energy_Bin_341  <= s_Energy_Bin_341  ;
  o_Energy_Bin_342  <= s_Energy_Bin_342  ;
  o_Energy_Bin_343  <= s_Energy_Bin_343  ;
  o_Energy_Bin_344  <= s_Energy_Bin_344  ;
  o_Energy_Bin_345  <= s_Energy_Bin_345  ;
  o_Energy_Bin_346  <= s_Energy_Bin_346  ;
  o_Energy_Bin_347  <= s_Energy_Bin_347  ;
  o_Energy_Bin_348  <= s_Energy_Bin_348  ;
  o_Energy_Bin_349  <= s_Energy_Bin_349  ;
  o_Energy_Bin_350  <= s_Energy_Bin_350  ;
  o_Energy_Bin_351  <= s_Energy_Bin_351  ;
  o_Energy_Bin_352  <= s_Energy_Bin_352  ;
  o_Energy_Bin_353  <= s_Energy_Bin_353  ;
  o_Energy_Bin_354  <= s_Energy_Bin_354  ;
  o_Energy_Bin_355  <= s_Energy_Bin_355  ;
  o_Energy_Bin_356  <= s_Energy_Bin_356  ;
  o_Energy_Bin_357  <= s_Energy_Bin_357  ;
  o_Energy_Bin_358  <= s_Energy_Bin_358  ;
  o_Energy_Bin_359  <= s_Energy_Bin_359  ;
  o_Energy_Bin_360  <= s_Energy_Bin_360  ;
  o_Energy_Bin_361  <= s_Energy_Bin_361  ;
  o_Energy_Bin_362  <= s_Energy_Bin_362  ;
  o_Energy_Bin_363  <= s_Energy_Bin_363  ;
  o_Energy_Bin_364  <= s_Energy_Bin_364  ;
  o_Energy_Bin_365  <= s_Energy_Bin_365  ;
  o_Energy_Bin_366  <= s_Energy_Bin_366  ;
  o_Energy_Bin_367  <= s_Energy_Bin_367  ;
  o_Energy_Bin_368  <= s_Energy_Bin_368  ;
  o_Energy_Bin_369  <= s_Energy_Bin_369  ;
  o_Energy_Bin_370  <= s_Energy_Bin_370  ;
  o_Energy_Bin_371  <= s_Energy_Bin_371  ;
  o_Energy_Bin_372  <= s_Energy_Bin_372  ;
  o_Energy_Bin_373  <= s_Energy_Bin_373  ;
  o_Energy_Bin_374  <= s_Energy_Bin_374  ;
  o_Energy_Bin_375  <= s_Energy_Bin_375  ;
  o_Energy_Bin_376  <= s_Energy_Bin_376  ;
  o_Energy_Bin_377  <= s_Energy_Bin_377  ;
  o_Energy_Bin_378  <= s_Energy_Bin_378  ;
  o_Energy_Bin_379  <= s_Energy_Bin_379  ;
  o_Energy_Bin_380  <= s_Energy_Bin_380  ;
  o_Energy_Bin_381  <= s_Energy_Bin_381  ;
  o_Energy_Bin_382  <= s_Energy_Bin_382  ;
  o_Energy_Bin_383  <= s_Energy_Bin_383  ;
  o_Energy_Bin_384  <= s_Energy_Bin_384  ;
  o_Energy_Bin_385  <= s_Energy_Bin_385  ;
  o_Energy_Bin_386  <= s_Energy_Bin_386  ;
  o_Energy_Bin_387  <= s_Energy_Bin_387  ;
  o_Energy_Bin_388  <= s_Energy_Bin_388  ;
  o_Energy_Bin_389  <= s_Energy_Bin_389  ;
  o_Energy_Bin_390  <= s_Energy_Bin_390  ;
  o_Energy_Bin_391  <= s_Energy_Bin_391  ;
  o_Energy_Bin_392  <= s_Energy_Bin_392  ;
  o_Energy_Bin_393  <= s_Energy_Bin_393  ;
  o_Energy_Bin_394  <= s_Energy_Bin_394  ;
  o_Energy_Bin_395  <= s_Energy_Bin_395  ;
  o_Energy_Bin_396  <= s_Energy_Bin_396  ;
  o_Energy_Bin_397  <= s_Energy_Bin_397  ;
  o_Energy_Bin_398  <= s_Energy_Bin_398  ;
  o_Energy_Bin_399  <= s_Energy_Bin_399  ;
  o_Energy_Bin_400  <= s_Energy_Bin_400  ;
  o_Energy_Bin_401  <= s_Energy_Bin_401  ;
  o_Energy_Bin_402  <= s_Energy_Bin_402  ;
  o_Energy_Bin_403  <= s_Energy_Bin_403  ;
  o_Energy_Bin_404  <= s_Energy_Bin_404  ;
  o_Energy_Bin_405  <= s_Energy_Bin_405  ;
  o_Energy_Bin_406  <= s_Energy_Bin_406  ;
  o_Energy_Bin_407  <= s_Energy_Bin_407  ;
  o_Energy_Bin_408  <= s_Energy_Bin_408  ;
  o_Energy_Bin_409  <= s_Energy_Bin_409  ;
  o_Energy_Bin_410  <= s_Energy_Bin_410  ;
  o_Energy_Bin_411  <= s_Energy_Bin_411  ;
  o_Energy_Bin_412  <= s_Energy_Bin_412  ;
  o_Energy_Bin_413  <= s_Energy_Bin_413  ;
  o_Energy_Bin_414  <= s_Energy_Bin_414  ;
  o_Energy_Bin_415  <= s_Energy_Bin_415  ;
  o_Energy_Bin_416  <= s_Energy_Bin_416  ;
  o_Energy_Bin_417  <= s_Energy_Bin_417  ;
  o_Energy_Bin_418  <= s_Energy_Bin_418  ;
  o_Energy_Bin_419  <= s_Energy_Bin_419  ;
  o_Energy_Bin_420  <= s_Energy_Bin_420  ;
  o_Energy_Bin_421  <= s_Energy_Bin_421  ;
  o_Energy_Bin_422  <= s_Energy_Bin_422  ;
  o_Energy_Bin_423  <= s_Energy_Bin_423  ;
  o_Energy_Bin_424  <= s_Energy_Bin_424  ;
  o_Energy_Bin_425  <= s_Energy_Bin_425  ;
  o_Energy_Bin_426  <= s_Energy_Bin_426  ;
  o_Energy_Bin_427  <= s_Energy_Bin_427  ;
  o_Energy_Bin_428  <= s_Energy_Bin_428  ;
  o_Energy_Bin_429  <= s_Energy_Bin_429  ;
  o_Energy_Bin_430  <= s_Energy_Bin_430  ;
  o_Energy_Bin_431  <= s_Energy_Bin_431  ;
  o_Energy_Bin_432  <= s_Energy_Bin_432  ;
  o_Energy_Bin_433  <= s_Energy_Bin_433  ;
  o_Energy_Bin_434  <= s_Energy_Bin_434  ;
  o_Energy_Bin_435  <= s_Energy_Bin_435  ;
  o_Energy_Bin_436  <= s_Energy_Bin_436  ;
  o_Energy_Bin_437  <= s_Energy_Bin_437  ;
  o_Energy_Bin_438  <= s_Energy_Bin_438  ;
  o_Energy_Bin_439  <= s_Energy_Bin_439  ;
  o_Energy_Bin_440  <= s_Energy_Bin_440  ;
  o_Energy_Bin_441  <= s_Energy_Bin_441  ;
  o_Energy_Bin_442  <= s_Energy_Bin_442  ;
  o_Energy_Bin_443  <= s_Energy_Bin_443  ;
  o_Energy_Bin_444  <= s_Energy_Bin_444  ;
  o_Energy_Bin_445  <= s_Energy_Bin_445  ;
  o_Energy_Bin_446  <= s_Energy_Bin_446  ;
  o_Energy_Bin_447  <= s_Energy_Bin_447  ;
  o_Energy_Bin_448  <= s_Energy_Bin_448  ;
  o_Energy_Bin_449  <= s_Energy_Bin_449  ;
  o_Energy_Bin_450  <= s_Energy_Bin_450  ;
  o_Energy_Bin_451  <= s_Energy_Bin_451  ;
  o_Energy_Bin_452  <= s_Energy_Bin_452  ;
  o_Energy_Bin_453  <= s_Energy_Bin_453  ;
  o_Energy_Bin_454  <= s_Energy_Bin_454  ;
  o_Energy_Bin_455  <= s_Energy_Bin_455  ;
  o_Energy_Bin_456  <= s_Energy_Bin_456  ;
  o_Energy_Bin_457  <= s_Energy_Bin_457  ;
  o_Energy_Bin_458  <= s_Energy_Bin_458  ;
  o_Energy_Bin_459  <= s_Energy_Bin_459  ;
  o_Energy_Bin_460  <= s_Energy_Bin_460  ;
  o_Energy_Bin_461  <= s_Energy_Bin_461  ;
  o_Energy_Bin_462  <= s_Energy_Bin_462  ;
  o_Energy_Bin_463  <= s_Energy_Bin_463  ;
  o_Energy_Bin_464  <= s_Energy_Bin_464  ;
  o_Energy_Bin_465  <= s_Energy_Bin_465  ;
  o_Energy_Bin_466  <= s_Energy_Bin_466  ;
  o_Energy_Bin_467  <= s_Energy_Bin_467  ;
  o_Energy_Bin_468  <= s_Energy_Bin_468  ;
  o_Energy_Bin_469  <= s_Energy_Bin_469  ;
  o_Energy_Bin_470  <= s_Energy_Bin_470  ;
  o_Energy_Bin_471  <= s_Energy_Bin_471  ;
  o_Energy_Bin_472  <= s_Energy_Bin_472  ;
  o_Energy_Bin_473  <= s_Energy_Bin_473  ;
  o_Energy_Bin_474  <= s_Energy_Bin_474  ;
  o_Energy_Bin_475  <= s_Energy_Bin_475  ;
  o_Energy_Bin_476  <= s_Energy_Bin_476  ;
  o_Energy_Bin_477  <= s_Energy_Bin_477  ;
  o_Energy_Bin_478  <= s_Energy_Bin_478  ;
  o_Energy_Bin_479  <= s_Energy_Bin_479  ;
  o_Energy_Bin_480  <= s_Energy_Bin_480  ;
  o_Energy_Bin_481  <= s_Energy_Bin_481  ;
  o_Energy_Bin_482  <= s_Energy_Bin_482  ;
  o_Energy_Bin_483  <= s_Energy_Bin_483  ;
  o_Energy_Bin_484  <= s_Energy_Bin_484  ;
  o_Energy_Bin_485  <= s_Energy_Bin_485  ;
  o_Energy_Bin_486  <= s_Energy_Bin_486  ;
  o_Energy_Bin_487  <= s_Energy_Bin_487  ;
  o_Energy_Bin_488  <= s_Energy_Bin_488  ;
  o_Energy_Bin_489  <= s_Energy_Bin_489  ;
  o_Energy_Bin_490  <= s_Energy_Bin_490  ;
  o_Energy_Bin_491  <= s_Energy_Bin_491  ;
  o_Energy_Bin_492  <= s_Energy_Bin_492  ;
  o_Energy_Bin_493  <= s_Energy_Bin_493  ;
  o_Energy_Bin_494  <= s_Energy_Bin_494  ;
  o_Energy_Bin_495  <= s_Energy_Bin_495  ;
  o_Energy_Bin_496  <= s_Energy_Bin_496  ;
  o_Energy_Bin_497  <= s_Energy_Bin_497  ;
  o_Energy_Bin_498  <= s_Energy_Bin_498  ;
  o_Energy_Bin_499  <= s_Energy_Bin_499  ;
  o_Energy_Bin_500  <= s_Energy_Bin_500  ;
  o_Energy_Bin_501  <= s_Energy_Bin_501  ;
  o_Energy_Bin_502  <= s_Energy_Bin_502  ;
  o_Energy_Bin_503  <= s_Energy_Bin_503  ;
  o_Energy_Bin_504  <= s_Energy_Bin_504  ;
  o_Energy_Bin_505  <= s_Energy_Bin_505  ;
  o_Energy_Bin_506  <= s_Energy_Bin_506  ;
  o_Energy_Bin_507  <= s_Energy_Bin_507  ;
  o_Energy_Bin_508  <= s_Energy_Bin_508  ;
  o_Energy_Bin_509  <= s_Energy_Bin_509  ;
  o_Energy_Bin_510  <= s_Energy_Bin_510  ;
  o_Energy_Bin_511  <= s_Energy_Bin_511  ;
  o_Energy_Bin_512  <= s_Energy_Bin_512  ;
  o_Energy_Bin_513  <= s_Energy_Bin_513  ;
  o_Energy_Bin_514  <= s_Energy_Bin_514  ;
  o_Energy_Bin_515  <= s_Energy_Bin_515  ;
  o_Energy_Bin_516  <= s_Energy_Bin_516  ;
  o_Energy_Bin_517  <= s_Energy_Bin_517  ;
  o_Energy_Bin_518  <= s_Energy_Bin_518  ;
  o_Energy_Bin_519  <= s_Energy_Bin_519  ;
  o_Energy_Bin_520  <= s_Energy_Bin_520  ;
  o_Energy_Bin_521  <= s_Energy_Bin_521  ;
  o_Energy_Bin_522  <= s_Energy_Bin_522  ;
  o_Energy_Bin_523  <= s_Energy_Bin_523  ;
  o_Energy_Bin_524  <= s_Energy_Bin_524  ;
  o_Energy_Bin_525  <= s_Energy_Bin_525  ;
  o_Energy_Bin_526  <= s_Energy_Bin_526  ;
  o_Energy_Bin_527  <= s_Energy_Bin_527  ;
  o_Energy_Bin_528  <= s_Energy_Bin_528  ;
  o_Energy_Bin_529  <= s_Energy_Bin_529  ;
  o_Energy_Bin_530  <= s_Energy_Bin_530  ;
  o_Energy_Bin_531  <= s_Energy_Bin_531  ;
  o_Energy_Bin_532  <= s_Energy_Bin_532  ;
  o_Energy_Bin_533  <= s_Energy_Bin_533  ;
  o_Energy_Bin_534  <= s_Energy_Bin_534  ;
  o_Energy_Bin_535  <= s_Energy_Bin_535  ;
  o_Energy_Bin_536  <= s_Energy_Bin_536  ;
  o_Energy_Bin_537  <= s_Energy_Bin_537  ;
  o_Energy_Bin_538  <= s_Energy_Bin_538  ;
  o_Energy_Bin_539  <= s_Energy_Bin_539  ;
  o_Energy_Bin_540  <= s_Energy_Bin_540  ;
  o_Energy_Bin_541  <= s_Energy_Bin_541  ;
  o_Energy_Bin_542  <= s_Energy_Bin_542  ;
  o_Energy_Bin_543  <= s_Energy_Bin_543  ;
  o_Energy_Bin_544  <= s_Energy_Bin_544  ;
  o_Energy_Bin_545  <= s_Energy_Bin_545  ;
  o_Energy_Bin_546  <= s_Energy_Bin_546  ;
  o_Energy_Bin_547  <= s_Energy_Bin_547  ;
  o_Energy_Bin_548  <= s_Energy_Bin_548  ;
  o_Energy_Bin_549  <= s_Energy_Bin_549  ;
  o_Energy_Bin_550  <= s_Energy_Bin_550  ;
  o_Energy_Bin_551  <= s_Energy_Bin_551  ;
  o_Energy_Bin_552  <= s_Energy_Bin_552  ;
  o_Energy_Bin_553  <= s_Energy_Bin_553  ;
  o_Energy_Bin_554  <= s_Energy_Bin_554  ;
  o_Energy_Bin_555  <= s_Energy_Bin_555  ;
  o_Energy_Bin_556  <= s_Energy_Bin_556  ;
  o_Energy_Bin_557  <= s_Energy_Bin_557  ;
  o_Energy_Bin_558  <= s_Energy_Bin_558  ;
  o_Energy_Bin_559  <= s_Energy_Bin_559  ;
  o_Energy_Bin_560  <= s_Energy_Bin_560  ;
  o_Energy_Bin_561  <= s_Energy_Bin_561  ;
  o_Energy_Bin_562  <= s_Energy_Bin_562  ;
  o_Energy_Bin_563  <= s_Energy_Bin_563  ;
  o_Energy_Bin_564  <= s_Energy_Bin_564  ;
  o_Energy_Bin_565  <= s_Energy_Bin_565  ;
  o_Energy_Bin_566  <= s_Energy_Bin_566  ;
  o_Energy_Bin_567  <= s_Energy_Bin_567  ;
  o_Energy_Bin_568  <= s_Energy_Bin_568  ;
  o_Energy_Bin_569  <= s_Energy_Bin_569  ;
  o_Energy_Bin_570  <= s_Energy_Bin_570  ;
  o_Energy_Bin_571  <= s_Energy_Bin_571  ;
  o_Energy_Bin_572  <= s_Energy_Bin_572  ;
  o_Energy_Bin_573  <= s_Energy_Bin_573  ;
  o_Energy_Bin_574  <= s_Energy_Bin_574  ;
  o_Energy_Bin_575  <= s_Energy_Bin_575  ;
  o_Energy_Bin_576  <= s_Energy_Bin_576  ;
  o_Energy_Bin_577  <= s_Energy_Bin_577  ;
  o_Energy_Bin_578  <= s_Energy_Bin_578  ;
  o_Energy_Bin_579  <= s_Energy_Bin_579  ;
  o_Energy_Bin_580  <= s_Energy_Bin_580  ;
  o_Energy_Bin_581  <= s_Energy_Bin_581  ;
  o_Energy_Bin_582  <= s_Energy_Bin_582  ;
  o_Energy_Bin_583  <= s_Energy_Bin_583  ;
  o_Energy_Bin_584  <= s_Energy_Bin_584  ;
  o_Energy_Bin_585  <= s_Energy_Bin_585  ;
  o_Energy_Bin_586  <= s_Energy_Bin_586  ;
  o_Energy_Bin_587  <= s_Energy_Bin_587  ;
  o_Energy_Bin_588  <= s_Energy_Bin_588  ;
  o_Energy_Bin_589  <= s_Energy_Bin_589  ;
  o_Energy_Bin_590  <= s_Energy_Bin_590  ;
  o_Energy_Bin_591  <= s_Energy_Bin_591  ;
  o_Energy_Bin_592  <= s_Energy_Bin_592  ;
  o_Energy_Bin_593  <= s_Energy_Bin_593  ;
  o_Energy_Bin_594  <= s_Energy_Bin_594  ;
  o_Energy_Bin_595  <= s_Energy_Bin_595  ;
  o_Energy_Bin_596  <= s_Energy_Bin_596  ;
  o_Energy_Bin_597  <= s_Energy_Bin_597  ;
  o_Energy_Bin_598  <= s_Energy_Bin_598  ;
  o_Energy_Bin_599  <= s_Energy_Bin_599  ;
  o_Energy_Bin_600  <= s_Energy_Bin_600  ;
  o_Energy_Bin_601  <= s_Energy_Bin_601  ;
  o_Energy_Bin_602  <= s_Energy_Bin_602  ;
  o_Energy_Bin_603  <= s_Energy_Bin_603  ;
  o_Energy_Bin_604  <= s_Energy_Bin_604  ;
  o_Energy_Bin_605  <= s_Energy_Bin_605  ;
  o_Energy_Bin_606  <= s_Energy_Bin_606  ;
  o_Energy_Bin_607  <= s_Energy_Bin_607  ;
  o_Energy_Bin_608  <= s_Energy_Bin_608  ;
  o_Energy_Bin_609  <= s_Energy_Bin_609  ;
  o_Energy_Bin_610  <= s_Energy_Bin_610  ;
  o_Energy_Bin_611  <= s_Energy_Bin_611  ;
  o_Energy_Bin_612  <= s_Energy_Bin_612  ;
  o_Energy_Bin_613  <= s_Energy_Bin_613  ;
  o_Energy_Bin_614  <= s_Energy_Bin_614  ;
  o_Energy_Bin_615  <= s_Energy_Bin_615  ;
  o_Energy_Bin_616  <= s_Energy_Bin_616  ;
  o_Energy_Bin_617  <= s_Energy_Bin_617  ;
  o_Energy_Bin_618  <= s_Energy_Bin_618  ;
  o_Energy_Bin_619  <= s_Energy_Bin_619  ;
  o_Energy_Bin_620  <= s_Energy_Bin_620  ;
  o_Energy_Bin_621  <= s_Energy_Bin_621  ;
  o_Energy_Bin_622  <= s_Energy_Bin_622  ;
  o_Energy_Bin_623  <= s_Energy_Bin_623  ;
  o_Energy_Bin_624  <= s_Energy_Bin_624  ;
  o_Energy_Bin_625  <= s_Energy_Bin_625  ;
  o_Energy_Bin_626  <= s_Energy_Bin_626  ;
  o_Energy_Bin_627  <= s_Energy_Bin_627  ;
  o_Energy_Bin_628  <= s_Energy_Bin_628  ;
  o_Energy_Bin_629  <= s_Energy_Bin_629  ;
  o_Energy_Bin_630  <= s_Energy_Bin_630  ;
  o_Energy_Bin_631  <= s_Energy_Bin_631  ;
  o_Energy_Bin_632  <= s_Energy_Bin_632  ;
  o_Energy_Bin_633  <= s_Energy_Bin_633  ;
  o_Energy_Bin_634  <= s_Energy_Bin_634  ;
  o_Energy_Bin_635  <= s_Energy_Bin_635  ;
  o_Energy_Bin_636  <= s_Energy_Bin_636  ;
  o_Energy_Bin_637  <= s_Energy_Bin_637  ;
  o_Energy_Bin_638  <= s_Energy_Bin_638  ;
  o_Energy_Bin_639  <= s_Energy_Bin_639  ;
  o_Energy_Bin_640  <= s_Energy_Bin_640  ;
  o_Energy_Bin_641  <= s_Energy_Bin_641  ;
  o_Energy_Bin_642  <= s_Energy_Bin_642  ;
  o_Energy_Bin_643  <= s_Energy_Bin_643  ;
  o_Energy_Bin_644  <= s_Energy_Bin_644  ;
  o_Energy_Bin_645  <= s_Energy_Bin_645  ;
  o_Energy_Bin_646  <= s_Energy_Bin_646  ;
  o_Energy_Bin_647  <= s_Energy_Bin_647  ;
  o_Energy_Bin_648  <= s_Energy_Bin_648  ;
  o_Energy_Bin_649  <= s_Energy_Bin_649  ;
  o_Energy_Bin_650  <= s_Energy_Bin_650  ;
  o_Energy_Bin_651  <= s_Energy_Bin_651  ;
  o_Energy_Bin_652  <= s_Energy_Bin_652  ;
  o_Energy_Bin_653  <= s_Energy_Bin_653  ;
  o_Energy_Bin_654  <= s_Energy_Bin_654  ;
  o_Energy_Bin_655  <= s_Energy_Bin_655  ;
  o_Energy_Bin_656  <= s_Energy_Bin_656  ;
  o_Energy_Bin_657  <= s_Energy_Bin_657  ;
  o_Energy_Bin_658  <= s_Energy_Bin_658  ;
  o_Energy_Bin_659  <= s_Energy_Bin_659  ;
  o_Energy_Bin_660  <= s_Energy_Bin_660  ;
  o_Energy_Bin_661  <= s_Energy_Bin_661  ;
  o_Energy_Bin_662  <= s_Energy_Bin_662  ;
  o_Energy_Bin_663  <= s_Energy_Bin_663  ;
  o_Energy_Bin_664  <= s_Energy_Bin_664  ;
  o_Energy_Bin_665  <= s_Energy_Bin_665  ;
  o_Energy_Bin_666  <= s_Energy_Bin_666  ;
  o_Energy_Bin_667  <= s_Energy_Bin_667  ;
  o_Energy_Bin_668  <= s_Energy_Bin_668  ;
  o_Energy_Bin_669  <= s_Energy_Bin_669  ;
  o_Energy_Bin_670  <= s_Energy_Bin_670  ;
  o_Energy_Bin_671  <= s_Energy_Bin_671  ;
  o_Energy_Bin_672  <= s_Energy_Bin_672  ;
  o_Energy_Bin_673  <= s_Energy_Bin_673  ;
  o_Energy_Bin_674  <= s_Energy_Bin_674  ;
  o_Energy_Bin_675  <= s_Energy_Bin_675  ;
  o_Energy_Bin_676  <= s_Energy_Bin_676  ;
  o_Energy_Bin_677  <= s_Energy_Bin_677  ;
  o_Energy_Bin_678  <= s_Energy_Bin_678  ;
  o_Energy_Bin_679  <= s_Energy_Bin_679  ;
  o_Energy_Bin_680  <= s_Energy_Bin_680  ;
  o_Energy_Bin_681  <= s_Energy_Bin_681  ;
  o_Energy_Bin_682  <= s_Energy_Bin_682  ;
  o_Energy_Bin_683  <= s_Energy_Bin_683  ;
  o_Energy_Bin_684  <= s_Energy_Bin_684  ;
  o_Energy_Bin_685  <= s_Energy_Bin_685  ;
  o_Energy_Bin_686  <= s_Energy_Bin_686  ;
  o_Energy_Bin_687  <= s_Energy_Bin_687  ;
  o_Energy_Bin_688  <= s_Energy_Bin_688  ;
  o_Energy_Bin_689  <= s_Energy_Bin_689  ;
  o_Energy_Bin_690  <= s_Energy_Bin_690  ;
  o_Energy_Bin_691  <= s_Energy_Bin_691  ;
  o_Energy_Bin_692  <= s_Energy_Bin_692  ;
  o_Energy_Bin_693  <= s_Energy_Bin_693  ;
  o_Energy_Bin_694  <= s_Energy_Bin_694  ;
  o_Energy_Bin_695  <= s_Energy_Bin_695  ;
  o_Energy_Bin_696  <= s_Energy_Bin_696  ;
  o_Energy_Bin_697  <= s_Energy_Bin_697  ;
  o_Energy_Bin_698  <= s_Energy_Bin_698  ;
  o_Energy_Bin_699  <= s_Energy_Bin_699  ;
  o_Energy_Bin_700  <= s_Energy_Bin_700  ;
  o_Energy_Bin_701  <= s_Energy_Bin_701  ;
  o_Energy_Bin_702  <= s_Energy_Bin_702  ;
  o_Energy_Bin_703  <= s_Energy_Bin_703  ;
  o_Energy_Bin_704  <= s_Energy_Bin_704  ;
  o_Energy_Bin_705  <= s_Energy_Bin_705  ;
  o_Energy_Bin_706  <= s_Energy_Bin_706  ;
  o_Energy_Bin_707  <= s_Energy_Bin_707  ;
  o_Energy_Bin_708  <= s_Energy_Bin_708  ;
  o_Energy_Bin_709  <= s_Energy_Bin_709  ;
  o_Energy_Bin_710  <= s_Energy_Bin_710  ;
  o_Energy_Bin_711  <= s_Energy_Bin_711  ;
  o_Energy_Bin_712  <= s_Energy_Bin_712  ;
  o_Energy_Bin_713  <= s_Energy_Bin_713  ;
  o_Energy_Bin_714  <= s_Energy_Bin_714  ;
  o_Energy_Bin_715  <= s_Energy_Bin_715  ;
  o_Energy_Bin_716  <= s_Energy_Bin_716  ;
  o_Energy_Bin_717  <= s_Energy_Bin_717  ;
  o_Energy_Bin_718  <= s_Energy_Bin_718  ;
  o_Energy_Bin_719  <= s_Energy_Bin_719  ;
  o_Energy_Bin_720  <= s_Energy_Bin_720  ;
  o_Energy_Bin_721  <= s_Energy_Bin_721  ;
  o_Energy_Bin_722  <= s_Energy_Bin_722  ;
  o_Energy_Bin_723  <= s_Energy_Bin_723  ;
  o_Energy_Bin_724  <= s_Energy_Bin_724  ;
  o_Energy_Bin_725  <= s_Energy_Bin_725  ;
  o_Energy_Bin_726  <= s_Energy_Bin_726  ;
  o_Energy_Bin_727  <= s_Energy_Bin_727  ;
  o_Energy_Bin_728  <= s_Energy_Bin_728  ;
  o_Energy_Bin_729  <= s_Energy_Bin_729  ;
  o_Energy_Bin_730  <= s_Energy_Bin_730  ;
  o_Energy_Bin_731  <= s_Energy_Bin_731  ;
  o_Energy_Bin_732  <= s_Energy_Bin_732  ;
  o_Energy_Bin_733  <= s_Energy_Bin_733  ;
  o_Energy_Bin_734  <= s_Energy_Bin_734  ;
  o_Energy_Bin_735  <= s_Energy_Bin_735  ;
  o_Energy_Bin_736  <= s_Energy_Bin_736  ;
  o_Energy_Bin_737  <= s_Energy_Bin_737  ;
  o_Energy_Bin_738  <= s_Energy_Bin_738  ;
  o_Energy_Bin_739  <= s_Energy_Bin_739  ;
  o_Energy_Bin_740  <= s_Energy_Bin_740  ;
  o_Energy_Bin_741  <= s_Energy_Bin_741  ;
  o_Energy_Bin_742  <= s_Energy_Bin_742  ;
  o_Energy_Bin_743  <= s_Energy_Bin_743  ;
  o_Energy_Bin_744  <= s_Energy_Bin_744  ;
  o_Energy_Bin_745  <= s_Energy_Bin_745  ;
  o_Energy_Bin_746  <= s_Energy_Bin_746  ;
  o_Energy_Bin_747  <= s_Energy_Bin_747  ;
  o_Energy_Bin_748  <= s_Energy_Bin_748  ;
  o_Energy_Bin_749  <= s_Energy_Bin_749  ;
  o_Energy_Bin_750  <= s_Energy_Bin_750  ;
  o_Energy_Bin_751  <= s_Energy_Bin_751  ;
  o_Energy_Bin_752  <= s_Energy_Bin_752  ;
  o_Energy_Bin_753  <= s_Energy_Bin_753  ;
  o_Energy_Bin_754  <= s_Energy_Bin_754  ;
  o_Energy_Bin_755  <= s_Energy_Bin_755  ;
  o_Energy_Bin_756  <= s_Energy_Bin_756  ;
  o_Energy_Bin_757  <= s_Energy_Bin_757  ;
  o_Energy_Bin_758  <= s_Energy_Bin_758  ;
  o_Energy_Bin_759  <= s_Energy_Bin_759  ;
  o_Energy_Bin_760  <= s_Energy_Bin_760  ;
  o_Energy_Bin_761  <= s_Energy_Bin_761  ;
  o_Energy_Bin_762  <= s_Energy_Bin_762  ;
  o_Energy_Bin_763  <= s_Energy_Bin_763  ;
  o_Energy_Bin_764  <= s_Energy_Bin_764  ;
  o_Energy_Bin_765  <= s_Energy_Bin_765  ;
  o_Energy_Bin_766  <= s_Energy_Bin_766  ;
  o_Energy_Bin_767  <= s_Energy_Bin_767  ;
  o_Energy_Bin_768  <= s_Energy_Bin_768  ;
  o_Energy_Bin_769  <= s_Energy_Bin_769  ;
  o_Energy_Bin_770  <= s_Energy_Bin_770  ;
  o_Energy_Bin_771  <= s_Energy_Bin_771  ;
  o_Energy_Bin_772  <= s_Energy_Bin_772  ;
  o_Energy_Bin_773  <= s_Energy_Bin_773  ;
  o_Energy_Bin_774  <= s_Energy_Bin_774  ;
  o_Energy_Bin_775  <= s_Energy_Bin_775  ;
  o_Energy_Bin_776  <= s_Energy_Bin_776  ;
  o_Energy_Bin_777  <= s_Energy_Bin_777  ;
  o_Energy_Bin_778  <= s_Energy_Bin_778  ;
  o_Energy_Bin_779  <= s_Energy_Bin_779  ;
  o_Energy_Bin_780  <= s_Energy_Bin_780  ;
  o_Energy_Bin_781  <= s_Energy_Bin_781  ;
  o_Energy_Bin_782  <= s_Energy_Bin_782  ;
  o_Energy_Bin_783  <= s_Energy_Bin_783  ;
  o_Energy_Bin_784  <= s_Energy_Bin_784  ;
  o_Energy_Bin_785  <= s_Energy_Bin_785  ;
  o_Energy_Bin_786  <= s_Energy_Bin_786  ;
  o_Energy_Bin_787  <= s_Energy_Bin_787  ;
  o_Energy_Bin_788  <= s_Energy_Bin_788  ;
  o_Energy_Bin_789  <= s_Energy_Bin_789  ;
  o_Energy_Bin_790  <= s_Energy_Bin_790  ;
  o_Energy_Bin_791  <= s_Energy_Bin_791  ;
  o_Energy_Bin_792  <= s_Energy_Bin_792  ;
  o_Energy_Bin_793  <= s_Energy_Bin_793  ;
  o_Energy_Bin_794  <= s_Energy_Bin_794  ;
  o_Energy_Bin_795  <= s_Energy_Bin_795  ;
  o_Energy_Bin_796  <= s_Energy_Bin_796  ;
  o_Energy_Bin_797  <= s_Energy_Bin_797  ;
  o_Energy_Bin_798  <= s_Energy_Bin_798  ;
  o_Energy_Bin_799  <= s_Energy_Bin_799  ;
  o_Energy_Bin_800  <= s_Energy_Bin_800  ;
  o_Energy_Bin_801  <= s_Energy_Bin_801  ;
  o_Energy_Bin_802  <= s_Energy_Bin_802  ;
  o_Energy_Bin_803  <= s_Energy_Bin_803  ;
  o_Energy_Bin_804  <= s_Energy_Bin_804  ;
  o_Energy_Bin_805  <= s_Energy_Bin_805  ;
  o_Energy_Bin_806  <= s_Energy_Bin_806  ;
  o_Energy_Bin_807  <= s_Energy_Bin_807  ;
  o_Energy_Bin_808  <= s_Energy_Bin_808  ;
  o_Energy_Bin_809  <= s_Energy_Bin_809  ;
  o_Energy_Bin_810  <= s_Energy_Bin_810  ;
  o_Energy_Bin_811  <= s_Energy_Bin_811  ;
  o_Energy_Bin_812  <= s_Energy_Bin_812  ;
  o_Energy_Bin_813  <= s_Energy_Bin_813  ;
  o_Energy_Bin_814  <= s_Energy_Bin_814  ;
  o_Energy_Bin_815  <= s_Energy_Bin_815  ;
  o_Energy_Bin_816  <= s_Energy_Bin_816  ;
  o_Energy_Bin_817  <= s_Energy_Bin_817  ;
  o_Energy_Bin_818  <= s_Energy_Bin_818  ;
  o_Energy_Bin_819  <= s_Energy_Bin_819  ;
  o_Energy_Bin_820  <= s_Energy_Bin_820  ;
  o_Energy_Bin_821  <= s_Energy_Bin_821  ;
  o_Energy_Bin_822  <= s_Energy_Bin_822  ;
  o_Energy_Bin_823  <= s_Energy_Bin_823  ;
  o_Energy_Bin_824  <= s_Energy_Bin_824  ;
  o_Energy_Bin_825  <= s_Energy_Bin_825  ;
  o_Energy_Bin_826  <= s_Energy_Bin_826  ;
  o_Energy_Bin_827  <= s_Energy_Bin_827  ;
  o_Energy_Bin_828  <= s_Energy_Bin_828  ;
  o_Energy_Bin_829  <= s_Energy_Bin_829  ;
  o_Energy_Bin_830  <= s_Energy_Bin_830  ;
  o_Energy_Bin_831  <= s_Energy_Bin_831  ;
  o_Energy_Bin_832  <= s_Energy_Bin_832  ;
  o_Energy_Bin_833  <= s_Energy_Bin_833  ;
  o_Energy_Bin_834  <= s_Energy_Bin_834  ;
  o_Energy_Bin_835  <= s_Energy_Bin_835  ;
  o_Energy_Bin_836  <= s_Energy_Bin_836  ;
  o_Energy_Bin_837  <= s_Energy_Bin_837  ;
  o_Energy_Bin_838  <= s_Energy_Bin_838  ;
  o_Energy_Bin_839  <= s_Energy_Bin_839  ;
  o_Energy_Bin_840  <= s_Energy_Bin_840  ;
  o_Energy_Bin_841  <= s_Energy_Bin_841  ;
  o_Energy_Bin_842  <= s_Energy_Bin_842  ;
  o_Energy_Bin_843  <= s_Energy_Bin_843  ;
  o_Energy_Bin_844  <= s_Energy_Bin_844  ;
  o_Energy_Bin_845  <= s_Energy_Bin_845  ;
  o_Energy_Bin_846  <= s_Energy_Bin_846  ;
  o_Energy_Bin_847  <= s_Energy_Bin_847  ;
  o_Energy_Bin_848  <= s_Energy_Bin_848  ;
  o_Energy_Bin_849  <= s_Energy_Bin_849  ;
  o_Energy_Bin_850  <= s_Energy_Bin_850  ;
  o_Energy_Bin_851  <= s_Energy_Bin_851  ;
  o_Energy_Bin_852  <= s_Energy_Bin_852  ;
  o_Energy_Bin_853  <= s_Energy_Bin_853  ;
  o_Energy_Bin_854  <= s_Energy_Bin_854  ;
  o_Energy_Bin_855  <= s_Energy_Bin_855  ;
  o_Energy_Bin_856  <= s_Energy_Bin_856  ;
  o_Energy_Bin_857  <= s_Energy_Bin_857  ;
  o_Energy_Bin_858  <= s_Energy_Bin_858  ;
  o_Energy_Bin_859  <= s_Energy_Bin_859  ;
  o_Energy_Bin_860  <= s_Energy_Bin_860  ;
  o_Energy_Bin_861  <= s_Energy_Bin_861  ;
  o_Energy_Bin_862  <= s_Energy_Bin_862  ;
  o_Energy_Bin_863  <= s_Energy_Bin_863  ;
  o_Energy_Bin_864  <= s_Energy_Bin_864  ;
  o_Energy_Bin_865  <= s_Energy_Bin_865  ;
  o_Energy_Bin_866  <= s_Energy_Bin_866  ;
  o_Energy_Bin_867  <= s_Energy_Bin_867  ;
  o_Energy_Bin_868  <= s_Energy_Bin_868  ;
  o_Energy_Bin_869  <= s_Energy_Bin_869  ;
  o_Energy_Bin_870  <= s_Energy_Bin_870  ;
  o_Energy_Bin_871  <= s_Energy_Bin_871  ;
  o_Energy_Bin_872  <= s_Energy_Bin_872  ;
  o_Energy_Bin_873  <= s_Energy_Bin_873  ;
  o_Energy_Bin_874  <= s_Energy_Bin_874  ;
  o_Energy_Bin_875  <= s_Energy_Bin_875  ;
  o_Energy_Bin_876  <= s_Energy_Bin_876  ;
  o_Energy_Bin_877  <= s_Energy_Bin_877  ;
  o_Energy_Bin_878  <= s_Energy_Bin_878  ;
  o_Energy_Bin_879  <= s_Energy_Bin_879  ;
  o_Energy_Bin_880  <= s_Energy_Bin_880  ;
  o_Energy_Bin_881  <= s_Energy_Bin_881  ;
  o_Energy_Bin_882  <= s_Energy_Bin_882  ;
  o_Energy_Bin_883  <= s_Energy_Bin_883  ;
  o_Energy_Bin_884  <= s_Energy_Bin_884  ;
  o_Energy_Bin_885  <= s_Energy_Bin_885  ;
  o_Energy_Bin_886  <= s_Energy_Bin_886  ;
  o_Energy_Bin_887  <= s_Energy_Bin_887  ;
  o_Energy_Bin_888  <= s_Energy_Bin_888  ;
  o_Energy_Bin_889  <= s_Energy_Bin_889  ;
  o_Energy_Bin_890  <= s_Energy_Bin_890  ;
  o_Energy_Bin_891  <= s_Energy_Bin_891  ;
  o_Energy_Bin_892  <= s_Energy_Bin_892  ;
  o_Energy_Bin_893  <= s_Energy_Bin_893  ;
  o_Energy_Bin_894  <= s_Energy_Bin_894  ;
  o_Energy_Bin_895  <= s_Energy_Bin_895  ;
  o_Energy_Bin_896  <= s_Energy_Bin_896  ;
  o_Energy_Bin_897  <= s_Energy_Bin_897  ;
  o_Energy_Bin_898  <= s_Energy_Bin_898  ;
  o_Energy_Bin_899  <= s_Energy_Bin_899  ;
  o_Energy_Bin_900  <= s_Energy_Bin_900  ;
  o_Energy_Bin_901  <= s_Energy_Bin_901  ;
  o_Energy_Bin_902  <= s_Energy_Bin_902  ;
  o_Energy_Bin_903  <= s_Energy_Bin_903  ;
  o_Energy_Bin_904  <= s_Energy_Bin_904  ;
  o_Energy_Bin_905  <= s_Energy_Bin_905  ;
  o_Energy_Bin_906  <= s_Energy_Bin_906  ;
  o_Energy_Bin_907  <= s_Energy_Bin_907  ;
  o_Energy_Bin_908  <= s_Energy_Bin_908  ;
  o_Energy_Bin_909  <= s_Energy_Bin_909  ;
  o_Energy_Bin_910  <= s_Energy_Bin_910  ;
  o_Energy_Bin_911  <= s_Energy_Bin_911  ;
  o_Energy_Bin_912  <= s_Energy_Bin_912  ;
  o_Energy_Bin_913  <= s_Energy_Bin_913  ;
  o_Energy_Bin_914  <= s_Energy_Bin_914  ;
  o_Energy_Bin_915  <= s_Energy_Bin_915  ;
  o_Energy_Bin_916  <= s_Energy_Bin_916  ;
  o_Energy_Bin_917  <= s_Energy_Bin_917  ;
  o_Energy_Bin_918  <= s_Energy_Bin_918  ;
  o_Energy_Bin_919  <= s_Energy_Bin_919  ;
  o_Energy_Bin_920  <= s_Energy_Bin_920  ;
  o_Energy_Bin_921  <= s_Energy_Bin_921  ;
  o_Energy_Bin_922  <= s_Energy_Bin_922  ;
  o_Energy_Bin_923  <= s_Energy_Bin_923  ;
  o_Energy_Bin_924  <= s_Energy_Bin_924  ;
  o_Energy_Bin_925  <= s_Energy_Bin_925  ;
  o_Energy_Bin_926  <= s_Energy_Bin_926  ;
  o_Energy_Bin_927  <= s_Energy_Bin_927  ;
  o_Energy_Bin_928  <= s_Energy_Bin_928  ;
  o_Energy_Bin_929  <= s_Energy_Bin_929  ;
  o_Energy_Bin_930  <= s_Energy_Bin_930  ;
  o_Energy_Bin_931  <= s_Energy_Bin_931  ;
  o_Energy_Bin_932  <= s_Energy_Bin_932  ;
  o_Energy_Bin_933  <= s_Energy_Bin_933  ;
  o_Energy_Bin_934  <= s_Energy_Bin_934  ;
  o_Energy_Bin_935  <= s_Energy_Bin_935  ;
  o_Energy_Bin_936  <= s_Energy_Bin_936  ;
  o_Energy_Bin_937  <= s_Energy_Bin_937  ;
  o_Energy_Bin_938  <= s_Energy_Bin_938  ;
  o_Energy_Bin_939  <= s_Energy_Bin_939  ;
  o_Energy_Bin_940  <= s_Energy_Bin_940  ;
  o_Energy_Bin_941  <= s_Energy_Bin_941  ;
  o_Energy_Bin_942  <= s_Energy_Bin_942  ;
  o_Energy_Bin_943  <= s_Energy_Bin_943  ;
  o_Energy_Bin_944  <= s_Energy_Bin_944  ;
  o_Energy_Bin_945  <= s_Energy_Bin_945  ;
  o_Energy_Bin_946  <= s_Energy_Bin_946  ;
  o_Energy_Bin_947  <= s_Energy_Bin_947  ;
  o_Energy_Bin_948  <= s_Energy_Bin_948  ;
  o_Energy_Bin_949  <= s_Energy_Bin_949  ;
  o_Energy_Bin_950  <= s_Energy_Bin_950  ;
  o_Energy_Bin_951  <= s_Energy_Bin_951  ;
  o_Energy_Bin_952  <= s_Energy_Bin_952  ;
  o_Energy_Bin_953  <= s_Energy_Bin_953  ;
  o_Energy_Bin_954  <= s_Energy_Bin_954  ;
  o_Energy_Bin_955  <= s_Energy_Bin_955  ;
  o_Energy_Bin_956  <= s_Energy_Bin_956  ;
  o_Energy_Bin_957  <= s_Energy_Bin_957  ;
  o_Energy_Bin_958  <= s_Energy_Bin_958  ;
  o_Energy_Bin_959  <= s_Energy_Bin_959  ;
  o_Energy_Bin_960  <= s_Energy_Bin_960  ;
  o_Energy_Bin_961  <= s_Energy_Bin_961  ;
  o_Energy_Bin_962  <= s_Energy_Bin_962  ;
  o_Energy_Bin_963  <= s_Energy_Bin_963  ;
  o_Energy_Bin_964  <= s_Energy_Bin_964  ;
  o_Energy_Bin_965  <= s_Energy_Bin_965  ;
  o_Energy_Bin_966  <= s_Energy_Bin_966  ;
  o_Energy_Bin_967  <= s_Energy_Bin_967  ;
  o_Energy_Bin_968  <= s_Energy_Bin_968  ;
  o_Energy_Bin_969  <= s_Energy_Bin_969  ;
  o_Energy_Bin_970  <= s_Energy_Bin_970  ;
  o_Energy_Bin_971  <= s_Energy_Bin_971  ;
  o_Energy_Bin_972  <= s_Energy_Bin_972  ;
  o_Energy_Bin_973  <= s_Energy_Bin_973  ;
  o_Energy_Bin_974  <= s_Energy_Bin_974  ;
  o_Energy_Bin_975  <= s_Energy_Bin_975  ;
  o_Energy_Bin_976  <= s_Energy_Bin_976  ;
  o_Energy_Bin_977  <= s_Energy_Bin_977  ;
  o_Energy_Bin_978  <= s_Energy_Bin_978  ;
  o_Energy_Bin_979  <= s_Energy_Bin_979  ;
  o_Energy_Bin_980  <= s_Energy_Bin_980  ;
  o_Energy_Bin_981  <= s_Energy_Bin_981  ;
  o_Energy_Bin_982  <= s_Energy_Bin_982  ;
  o_Energy_Bin_983  <= s_Energy_Bin_983  ;
  o_Energy_Bin_984  <= s_Energy_Bin_984  ;
  o_Energy_Bin_985  <= s_Energy_Bin_985  ;
  o_Energy_Bin_986  <= s_Energy_Bin_986  ;
  o_Energy_Bin_987  <= s_Energy_Bin_987  ;
  o_Energy_Bin_988  <= s_Energy_Bin_988  ;
  o_Energy_Bin_989  <= s_Energy_Bin_989  ;
  o_Energy_Bin_990  <= s_Energy_Bin_990  ;
  o_Energy_Bin_991  <= s_Energy_Bin_991  ;
  o_Energy_Bin_992  <= s_Energy_Bin_992  ;
  o_Energy_Bin_993  <= s_Energy_Bin_993  ;
  o_Energy_Bin_994  <= s_Energy_Bin_994  ;
  o_Energy_Bin_995  <= s_Energy_Bin_995  ;
  o_Energy_Bin_996  <= s_Energy_Bin_996  ;
  o_Energy_Bin_997  <= s_Energy_Bin_997  ;
  o_Energy_Bin_998  <= s_Energy_Bin_998  ;
  o_Energy_Bin_999  <= s_Energy_Bin_999  ;
  o_Energy_Bin_1000 <= s_Energy_Bin_1000 ;
  o_Energy_Bin_1001 <= s_Energy_Bin_1001 ;
  o_Energy_Bin_1002 <= s_Energy_Bin_1002 ;
  o_Energy_Bin_1003 <= s_Energy_Bin_1003 ;
  o_Energy_Bin_1004 <= s_Energy_Bin_1004 ;
  o_Energy_Bin_1005 <= s_Energy_Bin_1005 ;
  o_Energy_Bin_1006 <= s_Energy_Bin_1006 ;
  o_Energy_Bin_1007 <= s_Energy_Bin_1007 ;
  o_Energy_Bin_1008 <= s_Energy_Bin_1008 ;
  o_Energy_Bin_1009 <= s_Energy_Bin_1009 ;
  o_Energy_Bin_1010 <= s_Energy_Bin_1010 ;
  o_Energy_Bin_1011 <= s_Energy_Bin_1011 ;
  o_Energy_Bin_1012 <= s_Energy_Bin_1012 ;
  o_Energy_Bin_1013 <= s_Energy_Bin_1013 ;
  o_Energy_Bin_1014 <= s_Energy_Bin_1014 ;
  o_Energy_Bin_1015 <= s_Energy_Bin_1015 ;
  o_Energy_Bin_1016 <= s_Energy_Bin_1016 ;
  o_Energy_Bin_1017 <= s_Energy_Bin_1017 ;
  o_Energy_Bin_1018 <= s_Energy_Bin_1018 ;
  o_Energy_Bin_1019 <= s_Energy_Bin_1019 ;
  o_Energy_Bin_1020 <= s_Energy_Bin_1020 ;
  o_Energy_Bin_1021 <= s_Energy_Bin_1021 ;
  o_Energy_Bin_1022 <= s_Energy_Bin_1022 ;
  o_Energy_Bin_1023 <= s_Energy_Bin_1023 ;
  o_Energy_Bin_1024 <= s_Energy_Bin_1024 ;

  s_PEAK_THD       <= i_PEAK_THD;
  s_PEAK_THD_pos   <= i_PEAK_THD_pos;
  
  o_DATA_OUT_C1    <= s_DATA_OUT_C1;
  o_DATA_OUT_C2    <= s_DATA_OUT_C2;

  Energy_Bin_Rdy    <= Energy_Bin_Rdy_1 or Energy_Bin_Rdy_2 or Energy_Bin_Rdy_3 or Energy_Bin_Rdy_4 or Energy_Bin_Rdy_5 or Energy_Bin_Rdy_6 or Energy_Bin_Rdy_7 or Energy_Bin_Rdy_8 or Energy_Bin_Rdy_9;
  Energy_Bin_Rdy_bk <= not Energy_Bin_Rdy;
  
  
  DataProc_C1 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
         Data0_s_C1 <= (others =>'0');
         Data1_s_C1 <= (others =>'0');
         Data2_s_C1 <= (others =>'0');
         Data3_s_C1 <= (others =>'0');
         Data4_s_C1 <= (others =>'0');
         Data5_s_C1 <= (others =>'0');
         Data6_s_C1 <= (others =>'0');
         Data7_s_C1 <= (others =>'0');
         Data8_s_C1 <= (others =>'0');
         Data9_s_C1 <= (others =>'0');
         
         Data10_s_C1 <= (others =>'0');
         Data11_s_C1 <= (others =>'0');
         Data12_s_C1 <= (others =>'0');
         Data13_s_C1 <= (others =>'0');
         Data14_s_C1 <= (others =>'0');
         Data15_s_C1 <= (others =>'0');
         Data16_s_C1 <= (others =>'0');
         Data17_s_C1 <= (others =>'0');
         Data18_s_C1 <= (others =>'0');
         Data19_s_C1 <= (others =>'0');
         Data20_s_C1 <= (others =>'0');
         Data21_s_C1 <= (others =>'0');
         Data22_s_C1 <= (others =>'0');
         Data23_s_C1 <= (others =>'0');
         Data24_s_C1 <= (others =>'0');
		 
      elsif(DATARDY1 = '1') then
         Data0_s_C1   <= DATA1;
         
         Data1_s_C1   <= Data0_s_C1;
         Data2_s_C1   <= Data1_s_C1;   
		 Data3_s_C1   <= Data2_s_C1;
		 Data4_s_C1   <= Data3_s_C1;
         Data5_s_C1   <= Data4_s_C1;
		 Data6_s_C1   <= Data5_s_C1;
		 Data7_s_C1   <= Data6_s_C1;
		 Data8_s_C1   <= Data7_s_C1;
         Data9_s_C1   <= Data8_s_C1;
         
         
		 Data10_s_C1  <= Data9_s_C1;
		 Data11_s_C1  <= Data10_s_C1;
         Data12_s_C1  <= Data11_s_C1;
         Data13_s_C1  <= Data12_s_C1;   
		 Data14_s_C1  <= Data13_s_C1;
		 Data15_s_C1  <= Data14_s_C1;
         Data16_s_C1  <= Data15_s_C1;
		 Data17_s_C1  <= Data16_s_C1;
		 Data18_s_C1  <= Data17_s_C1;
		 Data19_s_C1  <= Data18_s_C1;
         Data20_s_C1  <= Data19_s_C1;
		 Data21_s_C1  <= Data20_s_C1;
		 Data22_s_C1  <= Data21_s_C1;
		 Data23_s_C1  <= Data22_s_C1;
		 Data24_s_C1  <= Data23_s_C1;
 
      end if;
    end if;
  end process  DataProc_C1;  
  
  DataProc_C2 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
         Data0_s_C2 <= (others =>'0');
         Data1_s_C2 <= (others =>'0');
         Data2_s_C2 <= (others =>'0');
         Data3_s_C2 <= (others =>'0');
         Data4_s_C2 <= (others =>'0');
         Data5_s_C2 <= (others =>'0');
         Data6_s_C2 <= (others =>'0');
         Data7_s_C2 <= (others =>'0');
         Data8_s_C2 <= (others =>'0');
         Data9_s_C2 <= (others =>'0');
         
         Data10_s_C2 <= (others =>'0');
         Data11_s_C2 <= (others =>'0');
         Data12_s_C2 <= (others =>'0');
         Data13_s_C2 <= (others =>'0');
         Data14_s_C2 <= (others =>'0');
         Data15_s_C2 <= (others =>'0');
         Data16_s_C2 <= (others =>'0');
         Data17_s_C2 <= (others =>'0');
         Data18_s_C2 <= (others =>'0');
         Data19_s_C2 <= (others =>'0');
         Data20_s_C2 <= (others =>'0');
         Data21_s_C2 <= (others =>'0');
         Data22_s_C2 <= (others =>'0');
         Data23_s_C2 <= (others =>'0');
         Data24_s_C2 <= (others =>'0');

      elsif(DATARDY2 = '1') then
         Data0_s_C2   <= DATA2;
         
         Data1_s_C2   <= Data0_s_C2;
         Data2_s_C2   <= Data1_s_C2;   
		 Data3_s_C2   <= Data2_s_C2;
		 Data4_s_C2   <= Data3_s_C2;
         Data5_s_C2   <= Data4_s_C2;
		 Data6_s_C2   <= Data5_s_C2;
		 Data7_s_C2   <= Data6_s_C2;
		 Data8_s_C2   <= Data7_s_C2;
         Data9_s_C2   <= Data8_s_C2;
         
		 Data10_s_C2  <= Data9_s_C2;
		 Data11_s_C2  <= Data10_s_C2;
         Data12_s_C2  <= Data11_s_C2;
         Data13_s_C2  <= Data12_s_C2;   
		 Data14_s_C2  <= Data13_s_C2;
		 Data15_s_C2  <= Data14_s_C2;
         Data16_s_C2  <= Data15_s_C2;
		 Data17_s_C2  <= Data16_s_C2;
		 Data18_s_C2  <= Data17_s_C2;
		 Data19_s_C2  <= Data18_s_C2;
         Data20_s_C2  <= Data19_s_C2;
		 Data21_s_C2  <= Data20_s_C2;
		 Data22_s_C2  <= Data21_s_C2;
		 Data23_s_C2  <= Data22_s_C2;
		 Data24_s_C2  <= Data23_s_C2;
  
      end if;
    end if;
  end process  DataProc_C2;  
  

  Data_Flag_Proc : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
            s_DATA_OUT_C1  <= (others =>'0');
		    ADD_TIMP_FLAG  <= '0';	
		    Energy_Ris_Dis <= '0';
	  elsif(PEAK_FL_Ris = '1') then
		    s_DATA_OUT_C1          <= PEAK_C1;
			ADD_TIMP_FLAG          <= '1';
			Energy_Ris_Dis         <= '1';
	  else
		    ADD_TIMP_FLAG          <= '0';
		    Energy_Ris_Dis         <= '0';
	  end if;
    end if;
  end process  Data_Flag_Proc; 

  Data_Flag_Proc_Pos : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
            s_DATA_OUT_C2  <= (others =>'0');
		    ADD_TIMP_FLAG_pos  <= '0';	
		    Energy_Ris_Dis_pos <= '0';
	  elsif(PEAK_FL_Ris_pos = '1') then
			s_DATA_OUT_C2          <= PEAK_C1_pos;
			ADD_TIMP_FLAG_pos      <= '1';
			Energy_Ris_Dis_pos     <= '1';
	  else
		    ADD_TIMP_FLAG_pos      <= '0';
		    Energy_Ris_Dis_pos     <= '0';
	  end if;
    end if;
  end process  Data_Flag_Proc_Pos; 


  --+----------
  -- PeakProc:
  --       This module compares the data in three registers 
  --       If the middle register datum is greater than the 
  --       data in the two other registers and it is also
  --       greater than the threshold, latch the data and
  --       set the peak detect flag.
  --+----------
 PeakProc_C1 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        PEAK_FL_C1 <= '0';
        PEAK_C1    <=  (others =>'0');
         
      elsif( (Data15_s_C1 < s_PEAK_THD) and (Data9_s_C1 > Data10_s_C1) and (Data10_s_C1 > Data11_s_C1) and (Data11_s_C1 > Data12_s_C1) and (Data12_s_C1 < Data13_s_C1) and (Data13_s_C1 < Data14_s_C1) and (Data14_s_C1 < Data15_s_C1) ) then
             PEAK_FL_C1 <= '1';
             PEAK_C1    <= Data12_s_C1; 
      else
             PEAK_FL_C1 <= '0';
      end if; 
	  
    end if;
  end process  PeakProc_C1;  
  
  PEAK_FL_C1_Rising_Edge : process(CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        PEAK_FL_C1_s1 <= '0';  
        PEAK_FL_C1_s2 <= '0';
      else
        PEAK_FL_C1_s1 <= PEAK_FL_C1;
        PEAK_FL_C1_s2 <= PEAK_FL_C1_s1;
      end if;
    end if;
  end process  PEAK_FL_C1_Rising_Edge;  
  
  PEAK_FL_C1_Rising_Edge_det : process(CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        PEAK_FL_Ris <= '0';  
      elsif((PEAK_FL_C1_s1 and not PEAK_FL_C1_s2)= '1') then 
        PEAK_FL_Ris <= '1';
      else
        PEAK_FL_Ris <= '0';
      end if;
    end if;
  end process  PEAK_FL_C1_Rising_Edge_det;  
  
  PEAK_FL_C1_Rising_Edge_delay : process(CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        PEAK_FL_Ris_s <= '0';  
      elsif(PEAK_FL_Ris = '1') then 
        PEAK_FL_Ris_s <= '1';
      else
        PEAK_FL_Ris_s <= '0';
      end if;
    end if;
  end process  PEAK_FL_C1_Rising_Edge_delay;  

-- positive peak rising
 PeakProc_C1_Pos : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        PEAK_FL_C1_pos <= '0';
        PEAK_C1_pos    <=  (others =>'0');
         
      elsif( (Data15_s_C1 > s_PEAK_THD_pos) and (Data9_s_C1 < Data10_s_C1) and (Data10_s_C1 < Data11_s_C1) and (Data11_s_C1 < Data12_s_C1) and (Data12_s_C1 > Data13_s_C1) and (Data13_s_C1 > Data14_s_C1) and (Data14_s_C1 > Data15_s_C1) ) then
             PEAK_FL_C1_pos <= '1';
             PEAK_C1_pos    <= Data12_s_C1; 
      else
             PEAK_FL_C1_pos <= '0';
      end if; 
	  
    end if;
  end process  PeakProc_C1_Pos;  
  
  PEAK_FL_C1_POS_Rising_Edge : process(CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        PEAK_FL_C1_pos_s1 <= '0';  
        PEAK_FL_C1_pos_s2 <= '0';
      else
        PEAK_FL_C1_pos_s1 <= PEAK_FL_C1_pos;
        PEAK_FL_C1_pos_s2 <= PEAK_FL_C1_pos_s1;
      end if;
    end if;
  end process  PEAK_FL_C1_Pos_Rising_Edge;  
  
  PEAK_FL_C1_Pos_Rising_Edge_det : process(CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        PEAK_FL_Ris_pos <= '0';  
      elsif((PEAK_FL_C1_pos_s1 and not PEAK_FL_C1_pos_s2)= '1') then 
        PEAK_FL_Ris_pos <= '1';
      else
        PEAK_FL_Ris_pos <= '0';
      end if;
    end if;
  end process  PEAK_FL_C1_Pos_Rising_Edge_det;  
  
  PEAK_FL_C1_Rising_Edge_delay_Pos : process(CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        PEAK_FL_Ris_pos_s <= '0';  
      elsif(PEAK_FL_Ris_pos = '1') then 
        PEAK_FL_Ris_pos_s <= '1';
      else
        PEAK_FL_Ris_pos_s <= '0';
      end if;
    end if;
  end process  PEAK_FL_C1_Rising_Edge_delay_Pos;   
 
-- channel_1 positive energy bin
 Energy_Bin_Pos_1 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E1_C1_L_Pos and PEAK_C1_Pos <= s_E1_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1 <= s_Energy_Bin_Pos_1 +'1';
		 Energy_Bin_Pos_Rdy_1 <= '1';
		else
		 s_Energy_Bin_Pos_1 <= s_Energy_Bin_Pos_1;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1;   
  
  Energy_Bin_Pos_2 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_2   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_2 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E2_C1_L_Pos and PEAK_C1_Pos <= s_E2_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_2 <= s_Energy_Bin_Pos_2 +'1';
		 Energy_Bin_Pos_Rdy_2 <= '1';
		else
		 s_Energy_Bin_Pos_2 <= s_Energy_Bin_Pos_2;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_2 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_2;   
  
  Energy_Bin_Pos_3 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_3   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_3 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E3_C1_L_Pos and PEAK_C1_Pos <= s_E3_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_3 <= s_Energy_Bin_Pos_3 +'1';
		 Energy_Bin_Pos_Rdy_3 <= '1';
		else
		 s_Energy_Bin_Pos_3 <= s_Energy_Bin_Pos_3;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_3 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_3;   
  
  Energy_Bin_Pos_4 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_4   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_4 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E4_C1_L_Pos and PEAK_C1_Pos <= s_E4_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_4 <= s_Energy_Bin_Pos_4 +'1';
		 Energy_Bin_Pos_Rdy_4 <= '1';
		else
		 s_Energy_Bin_Pos_4 <= s_Energy_Bin_Pos_4;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_4 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_4;   
 
 
  Energy_Bin_Pos_5 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_5   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_5 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E5_C1_L_Pos and PEAK_C1_Pos <= s_E5_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_5 <= s_Energy_Bin_Pos_5 +'1';
		 Energy_Bin_Pos_Rdy_5 <= '1';
		else
		 s_Energy_Bin_Pos_5 <= s_Energy_Bin_Pos_5;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_5 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_5;  
 
  
  Energy_Bin_Pos_6 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_6   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_6 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E6_C1_L_Pos and PEAK_C1_Pos <= s_E6_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_6 <= s_Energy_Bin_Pos_6 +'1';
		 Energy_Bin_Pos_Rdy_6 <= '1';
		else
		 s_Energy_Bin_Pos_6 <= s_Energy_Bin_Pos_6;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_6 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_6;   
  
 Energy_Bin_Pos_7 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_7   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_7 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E7_C1_L_Pos and PEAK_C1_Pos <= s_E7_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_7 <= s_Energy_Bin_Pos_7 +'1';
		 Energy_Bin_Pos_Rdy_7 <= '1';
		else
		 s_Energy_Bin_Pos_7 <= s_Energy_Bin_Pos_7;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_7 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_7;   
  
  Energy_Bin_Pos_8 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_8   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_8 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E8_C1_L_Pos and PEAK_C1_Pos <= s_E8_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_8 <= s_Energy_Bin_Pos_8 +'1';
		 Energy_Bin_Pos_Rdy_8 <= '1';
		else
		 s_Energy_Bin_Pos_8 <= s_Energy_Bin_Pos_8;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_8 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_8;   
  
  Energy_Bin_Pos_9 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_9   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_9 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E9_C1_L_Pos and PEAK_C1_Pos <= s_E9_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_9 <= s_Energy_Bin_Pos_9 +'1';
		 Energy_Bin_Pos_Rdy_9 <= '1';
		else
		 s_Energy_Bin_Pos_9 <= s_Energy_Bin_Pos_9;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_9 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_9;   
  
  Energy_Bin_Pos_10 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_10   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_10 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E10_C1_L_Pos and PEAK_C1_Pos <= s_E10_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_10 <= s_Energy_Bin_Pos_10 +'1';
		 Energy_Bin_Pos_Rdy_10 <= '1';
		else
		 s_Energy_Bin_Pos_10 <= s_Energy_Bin_Pos_10;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_10 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_10;   
  
  Energy_Bin_Pos_11 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_11   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_11 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E11_C1_L_Pos and PEAK_C1_Pos <= s_E11_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_11 <= s_Energy_Bin_Pos_11 +'1';
		 Energy_Bin_Pos_Rdy_11 <= '1';
		else
		 s_Energy_Bin_Pos_11 <= s_Energy_Bin_Pos_11;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_11 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_11;   
  
    Energy_Bin_Pos_12 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_12   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_12 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E12_C1_L_Pos and PEAK_C1_Pos <= s_E12_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_12 <= s_Energy_Bin_Pos_12 +'1';
		 Energy_Bin_Pos_Rdy_12 <= '1';
		else
		 s_Energy_Bin_Pos_12 <= s_Energy_Bin_Pos_12;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_12 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_12;   

    Energy_Bin_Pos_13 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_13   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_13 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E13_C1_L_Pos and PEAK_C1_Pos <= s_E13_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_13 <= s_Energy_Bin_Pos_13 +'1';
		 Energy_Bin_Pos_Rdy_13 <= '1';
		else
		 s_Energy_Bin_Pos_13 <= s_Energy_Bin_Pos_13;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_13 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_13;   
  
     Energy_Bin_Pos_14 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_14   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_14 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E14_C1_L_Pos and PEAK_C1_Pos <= s_E14_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_14 <= s_Energy_Bin_Pos_14 +'1';
		 Energy_Bin_Pos_Rdy_14 <= '1';
		else
		 s_Energy_Bin_Pos_14 <= s_Energy_Bin_Pos_14;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_14 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_14;    
  
     Energy_Bin_Pos_15 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_15   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_15 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E15_C1_L_Pos and PEAK_C1_Pos <= s_E15_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_15 <= s_Energy_Bin_Pos_15 +'1';
		 Energy_Bin_Pos_Rdy_15 <= '1';
		else
		 s_Energy_Bin_Pos_15 <= s_Energy_Bin_Pos_15;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_15 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_15;      
  
     Energy_Bin_Pos_16 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_16   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_16 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E16_C1_L_Pos and PEAK_C1_Pos <= s_E16_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_16 <= s_Energy_Bin_Pos_16 +'1';
		 Energy_Bin_Pos_Rdy_16 <= '1';
		else
		 s_Energy_Bin_Pos_16 <= s_Energy_Bin_Pos_16;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_16 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_16;     
  
     Energy_Bin_Pos_17 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_17   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_17 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E17_C1_L_Pos and PEAK_C1_Pos <= s_E17_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_17 <= s_Energy_Bin_Pos_17 +'1';
		 Energy_Bin_Pos_Rdy_17 <= '1';
		else
		 s_Energy_Bin_Pos_17 <= s_Energy_Bin_Pos_17;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_17 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_17;     
  
     Energy_Bin_Pos_18 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_18   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_18 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E18_C1_L_Pos and PEAK_C1_Pos <= s_E18_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_18 <= s_Energy_Bin_Pos_18 +'1';
		 Energy_Bin_Pos_Rdy_18 <= '1';
		else
		 s_Energy_Bin_Pos_18 <= s_Energy_Bin_Pos_18;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_18 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_18;       
  
     Energy_Bin_Pos_19 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_19   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_19 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E19_C1_L_Pos and PEAK_C1_Pos <= s_E19_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_19 <= s_Energy_Bin_Pos_19 +'1';
		 Energy_Bin_Pos_Rdy_19 <= '1';
		else
		 s_Energy_Bin_Pos_19 <= s_Energy_Bin_Pos_19;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_19 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_19;     
  
      Energy_Bin_Pos_20 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_20   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_20 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E20_C1_L_Pos and PEAK_C1_Pos <= s_E20_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_20 <= s_Energy_Bin_Pos_20 +'1';
		 Energy_Bin_Pos_Rdy_20 <= '1';
		else
		 s_Energy_Bin_Pos_20 <= s_Energy_Bin_Pos_20;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_20 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_20;      
  
  Energy_Bin_Pos_21 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_21   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_21 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E21_C1_L_Pos and PEAK_C1_Pos <= s_E21_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_21 <= s_Energy_Bin_Pos_21 +'1';
		 Energy_Bin_Pos_Rdy_21 <= '1';
		else
		 s_Energy_Bin_Pos_21 <= s_Energy_Bin_Pos_21;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_21 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_21;   
  
    Energy_Bin_Pos_22 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_22   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_22 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E22_C1_L_Pos and PEAK_C1_Pos <= s_E22_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_22 <= s_Energy_Bin_Pos_22 +'1';
		 Energy_Bin_Pos_Rdy_22 <= '1';
		else
		 s_Energy_Bin_Pos_22 <= s_Energy_Bin_Pos_22;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_22 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_22;   

    Energy_Bin_Pos_23 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_23   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_23 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E23_C1_L_Pos and PEAK_C1_Pos <= s_E23_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_23 <= s_Energy_Bin_Pos_23 +'1';
		 Energy_Bin_Pos_Rdy_23 <= '1';
		else
		 s_Energy_Bin_Pos_23 <= s_Energy_Bin_Pos_23;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_23 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_23;   
  
     Energy_Bin_Pos_24 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_24   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_24 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E24_C1_L_Pos and PEAK_C1_Pos <= s_E24_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_24 <= s_Energy_Bin_Pos_24 +'1';
		 Energy_Bin_Pos_Rdy_24 <= '1';
		else
		 s_Energy_Bin_Pos_24 <= s_Energy_Bin_Pos_24;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_24 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_24;    
  
     Energy_Bin_Pos_25 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_25   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_25 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E25_C1_L_Pos and PEAK_C1_Pos <= s_E25_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_25 <= s_Energy_Bin_Pos_25 +'1';
		 Energy_Bin_Pos_Rdy_25 <= '1';
		else
		 s_Energy_Bin_Pos_25 <= s_Energy_Bin_Pos_25;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_25 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_25;      
  
     Energy_Bin_Pos_26 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_26   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_26 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E26_C1_L_Pos and PEAK_C1_Pos <= s_E26_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_26 <= s_Energy_Bin_Pos_26 +'1';
		 Energy_Bin_Pos_Rdy_26 <= '1';
		else
		 s_Energy_Bin_Pos_26 <= s_Energy_Bin_Pos_26;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_26 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_26;     
  
     Energy_Bin_Pos_27 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_27   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_27 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E27_C1_L_Pos and PEAK_C1_Pos <= s_E27_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_27 <= s_Energy_Bin_Pos_27 +'1';
		 Energy_Bin_Pos_Rdy_27 <= '1';
		else
		 s_Energy_Bin_Pos_27 <= s_Energy_Bin_Pos_27;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_27 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_27;     
  
     Energy_Bin_Pos_28 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_28   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_28 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E28_C1_L_Pos and PEAK_C1_Pos <= s_E28_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_28 <= s_Energy_Bin_Pos_28 +'1';
		 Energy_Bin_Pos_Rdy_28 <= '1';
		else
		 s_Energy_Bin_Pos_28 <= s_Energy_Bin_Pos_28;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_28 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_28;       
  
     Energy_Bin_Pos_29 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_29   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_29 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E29_C1_L_Pos and PEAK_C1_Pos <= s_E29_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_29 <= s_Energy_Bin_Pos_29 +'1';
		 Energy_Bin_Pos_Rdy_29 <= '1';
		else
		 s_Energy_Bin_Pos_29 <= s_Energy_Bin_Pos_29;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_29 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_29;   

  Energy_Bin_Pos_30 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_30   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_30 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E30_C1_L_Pos and PEAK_C1_Pos <= s_E30_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_30 <= s_Energy_Bin_Pos_30 +'1';
		 Energy_Bin_Pos_Rdy_30 <= '1';
		else
		 s_Energy_Bin_Pos_30 <= s_Energy_Bin_Pos_30;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_30 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_30;     
  
  Energy_Bin_Pos_31 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_31   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_31 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E31_C1_L_Pos and PEAK_C1_Pos <= s_E31_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_31 <= s_Energy_Bin_Pos_31 +'1';
		 Energy_Bin_Pos_Rdy_31 <= '1';
		else
		 s_Energy_Bin_Pos_31 <= s_Energy_Bin_Pos_31;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_31 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_31;   
  
    Energy_Bin_Pos_32 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_32   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_32 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E32_C1_L_Pos and PEAK_C1_Pos <= s_E32_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_32 <= s_Energy_Bin_Pos_32 +'1';
		 Energy_Bin_Pos_Rdy_32 <= '1';
		else
		 s_Energy_Bin_Pos_32 <= s_Energy_Bin_Pos_32;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_32 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_32;   

    Energy_Bin_Pos_33 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_33   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_33 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E33_C1_L_Pos and PEAK_C1_Pos <= s_E33_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_33 <= s_Energy_Bin_Pos_33 +'1';
		 Energy_Bin_Pos_Rdy_33 <= '1';
		else
		 s_Energy_Bin_Pos_33 <= s_Energy_Bin_Pos_33;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_33 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_33;   
  
     Energy_Bin_Pos_34 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_34   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_34 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E34_C1_L_Pos and PEAK_C1_Pos <= s_E34_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_34 <= s_Energy_Bin_Pos_34 +'1';
		 Energy_Bin_Pos_Rdy_34 <= '1';
		else
		 s_Energy_Bin_Pos_34 <= s_Energy_Bin_Pos_34;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_34 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_34;    
  
     Energy_Bin_Pos_35 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_35   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_35 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E35_C1_L_Pos and PEAK_C1_Pos <= s_E35_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_35 <= s_Energy_Bin_Pos_35 +'1';
		 Energy_Bin_Pos_Rdy_35 <= '1';
		else
		 s_Energy_Bin_Pos_35 <= s_Energy_Bin_Pos_35;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_35 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_35;      
  
     Energy_Bin_Pos_36 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_36   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_36 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E36_C1_L_Pos and PEAK_C1_Pos <= s_E36_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_36 <= s_Energy_Bin_Pos_36 +'1';
		 Energy_Bin_Pos_Rdy_36 <= '1';
		else
		 s_Energy_Bin_Pos_36 <= s_Energy_Bin_Pos_36;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_36 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_36;     
  
     Energy_Bin_Pos_37 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_37   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_37 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E37_C1_L_Pos and PEAK_C1_Pos <= s_E37_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_37 <= s_Energy_Bin_Pos_37 +'1';
		 Energy_Bin_Pos_Rdy_37 <= '1';
		else
		 s_Energy_Bin_Pos_37 <= s_Energy_Bin_Pos_37;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_37 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_37;     
  
     Energy_Bin_Pos_38 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_38   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_38 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E38_C1_L_Pos and PEAK_C1_Pos <= s_E38_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_38 <= s_Energy_Bin_Pos_38 +'1';
		 Energy_Bin_Pos_Rdy_38 <= '1';
		else
		 s_Energy_Bin_Pos_38 <= s_Energy_Bin_Pos_38;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_38 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_38;       
  
     Energy_Bin_Pos_39 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_39   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_39 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E39_C1_L_Pos and PEAK_C1_Pos <= s_E39_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_39 <= s_Energy_Bin_Pos_39 +'1';
		 Energy_Bin_Pos_Rdy_39 <= '1';
		else
		 s_Energy_Bin_Pos_39 <= s_Energy_Bin_Pos_39;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_39 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_39;       

  Energy_Bin_Pos_40 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_40   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_40 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E40_C1_L_Pos and PEAK_C1_Pos <= s_E40_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_40 <= s_Energy_Bin_Pos_40 +'1';
		 Energy_Bin_Pos_Rdy_40 <= '1';
		else
		 s_Energy_Bin_Pos_40 <= s_Energy_Bin_Pos_40;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_40 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_40;   
  
  Energy_Bin_Pos_41 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_41   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_41 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E41_C1_L_Pos and PEAK_C1_Pos <= s_E41_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_41 <= s_Energy_Bin_Pos_41 +'1';
		 Energy_Bin_Pos_Rdy_41 <= '1';
		else
		 s_Energy_Bin_Pos_41 <= s_Energy_Bin_Pos_41;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_41 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_41;   
  
    Energy_Bin_Pos_42 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_42   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_42 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E42_C1_L_Pos and PEAK_C1_Pos <= s_E42_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_42 <= s_Energy_Bin_Pos_42 +'1';
		 Energy_Bin_Pos_Rdy_42 <= '1';
		else
		 s_Energy_Bin_Pos_42 <= s_Energy_Bin_Pos_42;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_42 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_42;   

    Energy_Bin_Pos_43 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_43   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_43 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E43_C1_L_Pos and PEAK_C1_Pos <= s_E43_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_43 <= s_Energy_Bin_Pos_43 +'1';
		 Energy_Bin_Pos_Rdy_43 <= '1';
		else
		 s_Energy_Bin_Pos_43 <= s_Energy_Bin_Pos_43;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_43 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_43;   
  
     Energy_Bin_Pos_44 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_44   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_44 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E44_C1_L_Pos and PEAK_C1_Pos <= s_E44_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_44 <= s_Energy_Bin_Pos_44 +'1';
		 Energy_Bin_Pos_Rdy_44 <= '1';
		else
		 s_Energy_Bin_Pos_44 <= s_Energy_Bin_Pos_44;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_44 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_44;    
  
     Energy_Bin_Pos_45 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_45   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_45 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E45_C1_L_Pos and PEAK_C1_Pos <= s_E45_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_45 <= s_Energy_Bin_Pos_45 +'1';
		 Energy_Bin_Pos_Rdy_45 <= '1';
		else
		 s_Energy_Bin_Pos_45 <= s_Energy_Bin_Pos_45;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_45 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_45;      
  
     Energy_Bin_Pos_46 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_46   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_46 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E46_C1_L_Pos and PEAK_C1_Pos <= s_E46_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_46 <= s_Energy_Bin_Pos_46 +'1';
		 Energy_Bin_Pos_Rdy_46 <= '1';
		else
		 s_Energy_Bin_Pos_46 <= s_Energy_Bin_Pos_46;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_46 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_46;     
  
     Energy_Bin_Pos_47 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_47   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_47 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E47_C1_L_Pos and PEAK_C1_Pos <= s_E47_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_47 <= s_Energy_Bin_Pos_47 +'1';
		 Energy_Bin_Pos_Rdy_47 <= '1';
		else
		 s_Energy_Bin_Pos_47 <= s_Energy_Bin_Pos_47;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_47 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_47;     
  
     Energy_Bin_Pos_48 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_48   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_48 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E48_C1_L_Pos and PEAK_C1_Pos <= s_E48_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_48 <= s_Energy_Bin_Pos_48 +'1';
		 Energy_Bin_Pos_Rdy_48 <= '1';
		else
		 s_Energy_Bin_Pos_48 <= s_Energy_Bin_Pos_48;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_48 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_48;       
  
     Energy_Bin_Pos_49 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_49   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_49 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E49_C1_L_Pos and PEAK_C1_Pos <= s_E49_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_49 <= s_Energy_Bin_Pos_49 +'1';
		 Energy_Bin_Pos_Rdy_49 <= '1';
		else
		 s_Energy_Bin_Pos_49 <= s_Energy_Bin_Pos_49;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_49 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_49;        
 
  Energy_Bin_Pos_50 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_50   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_50 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E50_C1_L_Pos and PEAK_C1_Pos <= s_E50_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_50 <= s_Energy_Bin_Pos_50 +'1';
		 Energy_Bin_Pos_Rdy_50 <= '1';
		else
		 s_Energy_Bin_Pos_50 <= s_Energy_Bin_Pos_50;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_50 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_50;   
  
  Energy_Bin_Pos_51 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_51   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_51 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E51_C1_L_Pos and PEAK_C1_Pos <= s_E51_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_51 <= s_Energy_Bin_Pos_51 +'1';
		 Energy_Bin_Pos_Rdy_51 <= '1';
		else
		 s_Energy_Bin_Pos_51 <= s_Energy_Bin_Pos_51;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_51 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_51;   
  
    Energy_Bin_Pos_52 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_52   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_52 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E52_C1_L_Pos and PEAK_C1_Pos <= s_E52_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_52 <= s_Energy_Bin_Pos_52 +'1';
		 Energy_Bin_Pos_Rdy_52 <= '1';
		else
		 s_Energy_Bin_Pos_52 <= s_Energy_Bin_Pos_52;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_52 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_52;   

    Energy_Bin_Pos_53 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_53   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_53 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E53_C1_L_Pos and PEAK_C1_Pos <= s_E53_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_53 <= s_Energy_Bin_Pos_53 +'1';
		 Energy_Bin_Pos_Rdy_53 <= '1';
		else
		 s_Energy_Bin_Pos_53 <= s_Energy_Bin_Pos_53;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_53 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_53;   
  
     Energy_Bin_Pos_54 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_54   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_54 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E54_C1_L_Pos and PEAK_C1_Pos <= s_E54_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_54 <= s_Energy_Bin_Pos_54 +'1';
		 Energy_Bin_Pos_Rdy_54 <= '1';
		else
		 s_Energy_Bin_Pos_54 <= s_Energy_Bin_Pos_54;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_54 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_54;    
  
     Energy_Bin_Pos_55 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_55   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_55 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E55_C1_L_Pos and PEAK_C1_Pos <= s_E55_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_55 <= s_Energy_Bin_Pos_55 +'1';
		 Energy_Bin_Pos_Rdy_55 <= '1';
		else
		 s_Energy_Bin_Pos_55 <= s_Energy_Bin_Pos_55;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_55 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_55;      
  
     Energy_Bin_Pos_56 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_56   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_56 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E56_C1_L_Pos and PEAK_C1_Pos <= s_E56_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_56 <= s_Energy_Bin_Pos_56 +'1';
		 Energy_Bin_Pos_Rdy_56 <= '1';
		else
		 s_Energy_Bin_Pos_56 <= s_Energy_Bin_Pos_56;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_56 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_56;     
  
     Energy_Bin_Pos_57 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_57   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_57 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E57_C1_L_Pos and PEAK_C1_Pos <= s_E57_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_57 <= s_Energy_Bin_Pos_57 +'1';
		 Energy_Bin_Pos_Rdy_57 <= '1';
		else
		 s_Energy_Bin_Pos_57 <= s_Energy_Bin_Pos_57;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_57 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_57;     
  
     Energy_Bin_Pos_58 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_58   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_58 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E58_C1_L_Pos and PEAK_C1_Pos <= s_E58_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_58 <= s_Energy_Bin_Pos_58 +'1';
		 Energy_Bin_Pos_Rdy_58 <= '1';
		else
		 s_Energy_Bin_Pos_58 <= s_Energy_Bin_Pos_58;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_58 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_58;       
  
     Energy_Bin_Pos_59 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_59   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_59 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E59_C1_L_Pos and PEAK_C1_Pos <= s_E59_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_59 <= s_Energy_Bin_Pos_59 +'1';
		 Energy_Bin_Pos_Rdy_59 <= '1';
		else
		 s_Energy_Bin_Pos_59 <= s_Energy_Bin_Pos_59;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_59 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_59;        

     Energy_Bin_Pos_60 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_60   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_60 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E60_C1_L_Pos and PEAK_C1_Pos <= s_E60_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_60 <= s_Energy_Bin_Pos_60 +'1';
		 Energy_Bin_Pos_Rdy_60 <= '1';
		else
		 s_Energy_Bin_Pos_60 <= s_Energy_Bin_Pos_60;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_60 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_60; 
  
  Energy_Bin_Pos_61 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_61   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_61 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E61_C1_L_Pos and PEAK_C1_Pos <= s_E61_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_61 <= s_Energy_Bin_Pos_61 +'1';
		 Energy_Bin_Pos_Rdy_61 <= '1';
		else
		 s_Energy_Bin_Pos_61 <= s_Energy_Bin_Pos_61;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_61 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_61;   
  
    Energy_Bin_Pos_62 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_62   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_62 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E62_C1_L_Pos and PEAK_C1_Pos <= s_E62_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_62 <= s_Energy_Bin_Pos_62 +'1';
		 Energy_Bin_Pos_Rdy_62 <= '1';
		else
		 s_Energy_Bin_Pos_62 <= s_Energy_Bin_Pos_62;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_62 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_62;   

    Energy_Bin_Pos_63 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_63   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_63 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E63_C1_L_Pos and PEAK_C1_Pos <= s_E63_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_63 <= s_Energy_Bin_Pos_63 +'1';
		 Energy_Bin_Pos_Rdy_63 <= '1';
		else
		 s_Energy_Bin_Pos_63 <= s_Energy_Bin_Pos_63;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_63 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_63;   
  
     Energy_Bin_Pos_64 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_64   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_64 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E64_C1_L_Pos and PEAK_C1_Pos <= s_E64_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_64 <= s_Energy_Bin_Pos_64 +'1';
		 Energy_Bin_Pos_Rdy_64 <= '1';
		else
		 s_Energy_Bin_Pos_64 <= s_Energy_Bin_Pos_64;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_64 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_64;    
  
     Energy_Bin_Pos_65 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_65   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_65 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E65_C1_L_Pos and PEAK_C1_Pos <= s_E65_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_65 <= s_Energy_Bin_Pos_65 +'1';
		 Energy_Bin_Pos_Rdy_65 <= '1';
		else
		 s_Energy_Bin_Pos_65 <= s_Energy_Bin_Pos_65;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_65 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_65;      
  
     Energy_Bin_Pos_66 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_66   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_66 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E66_C1_L_Pos and PEAK_C1_Pos <= s_E66_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_66 <= s_Energy_Bin_Pos_66 +'1';
		 Energy_Bin_Pos_Rdy_66 <= '1';
		else
		 s_Energy_Bin_Pos_66 <= s_Energy_Bin_Pos_66;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_66 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_66;     
  
     Energy_Bin_Pos_67 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_67   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_67 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E67_C1_L_Pos and PEAK_C1_Pos <= s_E67_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_67 <= s_Energy_Bin_Pos_67 +'1';
		 Energy_Bin_Pos_Rdy_67 <= '1';
		else
		 s_Energy_Bin_Pos_67 <= s_Energy_Bin_Pos_67;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_67 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_67;     
  
     Energy_Bin_Pos_68 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_68   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_68 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E68_C1_L_Pos and PEAK_C1_Pos <= s_E68_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_68 <= s_Energy_Bin_Pos_68 +'1';
		 Energy_Bin_Pos_Rdy_68 <= '1';
		else
		 s_Energy_Bin_Pos_68 <= s_Energy_Bin_Pos_68;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_68 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_68;       
  
     Energy_Bin_Pos_69 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_69   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_69 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E69_C1_L_Pos and PEAK_C1_Pos <= s_E69_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_69 <= s_Energy_Bin_Pos_69 +'1';
		 Energy_Bin_Pos_Rdy_69 <= '1';
		else
		 s_Energy_Bin_Pos_69 <= s_Energy_Bin_Pos_69;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_69 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_69;      

     Energy_Bin_Pos_70 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_70   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_70 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E70_C1_L_Pos and PEAK_C1_Pos <= s_E70_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_70 <= s_Energy_Bin_Pos_70 +'1';
		 Energy_Bin_Pos_Rdy_70 <= '1';
		else
		 s_Energy_Bin_Pos_70 <= s_Energy_Bin_Pos_70;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_70 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_70;       
  
  Energy_Bin_Pos_71 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_71   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_71 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E71_C1_L_Pos and PEAK_C1_Pos <= s_E71_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_71 <= s_Energy_Bin_Pos_71 +'1';
		 Energy_Bin_Pos_Rdy_71 <= '1';
		else
		 s_Energy_Bin_Pos_71 <= s_Energy_Bin_Pos_71;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_71 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_71;   
  
    Energy_Bin_Pos_72 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_72   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_72 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E72_C1_L_Pos and PEAK_C1_Pos <= s_E72_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_72 <= s_Energy_Bin_Pos_72 +'1';
		 Energy_Bin_Pos_Rdy_72 <= '1';
		else
		 s_Energy_Bin_Pos_72 <= s_Energy_Bin_Pos_72;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_72 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_72;   

    Energy_Bin_Pos_73 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_73   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_73 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E73_C1_L_Pos and PEAK_C1_Pos <= s_E73_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_73 <= s_Energy_Bin_Pos_73 +'1';
		 Energy_Bin_Pos_Rdy_73 <= '1';
		else
		 s_Energy_Bin_Pos_73 <= s_Energy_Bin_Pos_73;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_73 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_73;   
  
     Energy_Bin_Pos_74 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_74   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_74 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E74_C1_L_Pos and PEAK_C1_Pos <= s_E74_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_74 <= s_Energy_Bin_Pos_74 +'1';
		 Energy_Bin_Pos_Rdy_74 <= '1';
		else
		 s_Energy_Bin_Pos_74 <= s_Energy_Bin_Pos_74;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_74 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_74;    
  
     Energy_Bin_Pos_75 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_75   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_75 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E75_C1_L_Pos and PEAK_C1_Pos <= s_E75_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_75 <= s_Energy_Bin_Pos_75 +'1';
		 Energy_Bin_Pos_Rdy_75 <= '1';
		else
		 s_Energy_Bin_Pos_75 <= s_Energy_Bin_Pos_75;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_75 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_75;      
  
     Energy_Bin_Pos_76 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_76   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_76 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E76_C1_L_Pos and PEAK_C1_Pos <= s_E76_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_76 <= s_Energy_Bin_Pos_76 +'1';
		 Energy_Bin_Pos_Rdy_76 <= '1';
		else
		 s_Energy_Bin_Pos_76 <= s_Energy_Bin_Pos_76;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_76 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_76;     
  
     Energy_Bin_Pos_77 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_77   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_77 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E77_C1_L_Pos and PEAK_C1_Pos <= s_E77_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_77 <= s_Energy_Bin_Pos_77 +'1';
		 Energy_Bin_Pos_Rdy_77 <= '1';
		else
		 s_Energy_Bin_Pos_77 <= s_Energy_Bin_Pos_77;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_77 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_77;     
  
     Energy_Bin_Pos_78 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_78   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_78 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E78_C1_L_Pos and PEAK_C1_Pos <= s_E78_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_78 <= s_Energy_Bin_Pos_78 +'1';
		 Energy_Bin_Pos_Rdy_78 <= '1';
		else
		 s_Energy_Bin_Pos_78 <= s_Energy_Bin_Pos_78;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_78 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_78;       
  
     Energy_Bin_Pos_79 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_79   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_79 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E79_C1_L_Pos and PEAK_C1_Pos <= s_E79_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_79 <= s_Energy_Bin_Pos_79 +'1';
		 Energy_Bin_Pos_Rdy_79 <= '1';
		else
		 s_Energy_Bin_Pos_79 <= s_Energy_Bin_Pos_79;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_79 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_79;    
  
     Energy_Bin_Pos_80 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_80   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_80 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E80_C1_L_Pos and PEAK_C1_Pos <= s_E80_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_80 <= s_Energy_Bin_Pos_80 +'1';
		 Energy_Bin_Pos_Rdy_80 <= '1';
		else
		 s_Energy_Bin_Pos_80 <= s_Energy_Bin_Pos_80;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_80 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_80;       
  
  Energy_Bin_Pos_81 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_81   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_81 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E81_C1_L_Pos and PEAK_C1_Pos <= s_E81_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_81 <= s_Energy_Bin_Pos_81 +'1';
		 Energy_Bin_Pos_Rdy_81 <= '1';
		else
		 s_Energy_Bin_Pos_81 <= s_Energy_Bin_Pos_81;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_81 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_81;   
  
    Energy_Bin_Pos_82 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_82   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_82 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E82_C1_L_Pos and PEAK_C1_Pos <= s_E82_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_82 <= s_Energy_Bin_Pos_82 +'1';
		 Energy_Bin_Pos_Rdy_82 <= '1';
		else
		 s_Energy_Bin_Pos_82 <= s_Energy_Bin_Pos_82;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_82 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_82;   

    Energy_Bin_Pos_83 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_83   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_83 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E83_C1_L_Pos and PEAK_C1_Pos <= s_E83_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_83 <= s_Energy_Bin_Pos_83 +'1';
		 Energy_Bin_Pos_Rdy_83 <= '1';
		else
		 s_Energy_Bin_Pos_83 <= s_Energy_Bin_Pos_83;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_83 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_83;   
  
     Energy_Bin_Pos_84 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_84   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_84 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E84_C1_L_Pos and PEAK_C1_Pos <= s_E84_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_84 <= s_Energy_Bin_Pos_84 +'1';
		 Energy_Bin_Pos_Rdy_84 <= '1';
		else
		 s_Energy_Bin_Pos_84 <= s_Energy_Bin_Pos_84;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_84 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_84;    
  
     Energy_Bin_Pos_85 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_85   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_85 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E85_C1_L_Pos and PEAK_C1_Pos <= s_E85_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_85 <= s_Energy_Bin_Pos_85 +'1';
		 Energy_Bin_Pos_Rdy_85 <= '1';
		else
		 s_Energy_Bin_Pos_85 <= s_Energy_Bin_Pos_85;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_85 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_85;      
  
     Energy_Bin_Pos_86 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_86   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_86 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E86_C1_L_Pos and PEAK_C1_Pos <= s_E86_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_86 <= s_Energy_Bin_Pos_86 +'1';
		 Energy_Bin_Pos_Rdy_86 <= '1';
		else
		 s_Energy_Bin_Pos_86 <= s_Energy_Bin_Pos_86;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_86 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_86;     
  
     Energy_Bin_Pos_87 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_87   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_87 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E87_C1_L_Pos and PEAK_C1_Pos <= s_E87_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_87 <= s_Energy_Bin_Pos_87 +'1';
		 Energy_Bin_Pos_Rdy_87 <= '1';
		else
		 s_Energy_Bin_Pos_87 <= s_Energy_Bin_Pos_87;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_87 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_87;     
  
     Energy_Bin_Pos_88 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_88   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_88 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E88_C1_L_Pos and PEAK_C1_Pos <= s_E88_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_88 <= s_Energy_Bin_Pos_88 +'1';
		 Energy_Bin_Pos_Rdy_88 <= '1';
		else
		 s_Energy_Bin_Pos_88 <= s_Energy_Bin_Pos_88;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_88 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_88;       
  
     Energy_Bin_Pos_89 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_89   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_89 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E89_C1_L_Pos and PEAK_C1_Pos <= s_E89_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_89 <= s_Energy_Bin_Pos_89 +'1';
		 Energy_Bin_Pos_Rdy_89 <= '1';
		else
		 s_Energy_Bin_Pos_89 <= s_Energy_Bin_Pos_89;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_89 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_89;      

     Energy_Bin_Pos_90 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_90   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_90 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E90_C1_L_Pos and PEAK_C1_Pos <= s_E90_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_90 <= s_Energy_Bin_Pos_90 +'1';
		 Energy_Bin_Pos_Rdy_90 <= '1';
		else
		 s_Energy_Bin_Pos_90 <= s_Energy_Bin_Pos_90;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_90 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_90;       
  
  Energy_Bin_Pos_91 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_91   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_91 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E91_C1_L_Pos and PEAK_C1_Pos <= s_E91_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_91 <= s_Energy_Bin_Pos_91 +'1';
		 Energy_Bin_Pos_Rdy_91 <= '1';
		else
		 s_Energy_Bin_Pos_91 <= s_Energy_Bin_Pos_91;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_91 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_91;   
  
    Energy_Bin_Pos_92 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_92   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_92 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E92_C1_L_Pos and PEAK_C1_Pos <= s_E92_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_92 <= s_Energy_Bin_Pos_92 +'1';
		 Energy_Bin_Pos_Rdy_92 <= '1';
		else
		 s_Energy_Bin_Pos_92 <= s_Energy_Bin_Pos_92;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_92 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_92;   

    Energy_Bin_Pos_93 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_93   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_93 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E93_C1_L_Pos and PEAK_C1_Pos <= s_E93_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_93 <= s_Energy_Bin_Pos_93 +'1';
		 Energy_Bin_Pos_Rdy_93 <= '1';
		else
		 s_Energy_Bin_Pos_93 <= s_Energy_Bin_Pos_93;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_93 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_93;   
  
     Energy_Bin_Pos_94 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_94   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_94 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E94_C1_L_Pos and PEAK_C1_Pos <= s_E94_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_94 <= s_Energy_Bin_Pos_94 +'1';
		 Energy_Bin_Pos_Rdy_94 <= '1';
		else
		 s_Energy_Bin_Pos_94 <= s_Energy_Bin_Pos_94;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_94 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_94;    
  
     Energy_Bin_Pos_95 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_95   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_95 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E95_C1_L_Pos and PEAK_C1_Pos <= s_E95_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_95 <= s_Energy_Bin_Pos_95 +'1';
		 Energy_Bin_Pos_Rdy_95 <= '1';
		else
		 s_Energy_Bin_Pos_95 <= s_Energy_Bin_Pos_95;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_95 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_95;      
  
     Energy_Bin_Pos_96 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_96   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_96 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E96_C1_L_Pos and PEAK_C1_Pos <= s_E96_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_96 <= s_Energy_Bin_Pos_96 +'1';
		 Energy_Bin_Pos_Rdy_96 <= '1';
		else
		 s_Energy_Bin_Pos_96 <= s_Energy_Bin_Pos_96;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_96 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_96;     
  
     Energy_Bin_Pos_97 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_97   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_97 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E97_C1_L_Pos and PEAK_C1_Pos <= s_E97_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_97 <= s_Energy_Bin_Pos_97 +'1';
		 Energy_Bin_Pos_Rdy_97 <= '1';
		else
		 s_Energy_Bin_Pos_97 <= s_Energy_Bin_Pos_97;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_97 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_97;     
  
     Energy_Bin_Pos_98 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_98   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_98 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E98_C1_L_Pos and PEAK_C1_Pos <= s_E98_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_98 <= s_Energy_Bin_Pos_98 +'1';
		 Energy_Bin_Pos_Rdy_98 <= '1';
		else
		 s_Energy_Bin_Pos_98 <= s_Energy_Bin_Pos_98;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_98 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_98;       
  
     Energy_Bin_Pos_99 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_99   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_99 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E99_C1_L_Pos and PEAK_C1_Pos <= s_E99_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_99 <= s_Energy_Bin_Pos_99 +'1';
		 Energy_Bin_Pos_Rdy_99 <= '1';
		else
		 s_Energy_Bin_Pos_99 <= s_Energy_Bin_Pos_99;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_99 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_99;      
  
     Energy_Bin_Pos_100 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_100   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_100 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E100_C1_L_Pos and PEAK_C1_Pos <= s_E100_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_100 <= s_Energy_Bin_Pos_100 +'1';
		 Energy_Bin_Pos_Rdy_100 <= '1';
		else
		 s_Energy_Bin_Pos_100 <= s_Energy_Bin_Pos_100;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_100 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_100;    
  
  Energy_Bin_Pos_101 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_101   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_101 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E101_C1_L_Pos and PEAK_C1_Pos <= s_E101_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_101 <= s_Energy_Bin_Pos_101 +'1';
		 Energy_Bin_Pos_Rdy_101 <= '1';
		else
		 s_Energy_Bin_Pos_101 <= s_Energy_Bin_Pos_101;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_101 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_101;   
  
  Energy_Bin_Pos_102 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_102   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_102 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E102_C1_L_Pos and PEAK_C1_Pos <= s_E102_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_102 <= s_Energy_Bin_Pos_102 +'1';
		 Energy_Bin_Pos_Rdy_102 <= '1';
		else
		 s_Energy_Bin_Pos_102 <= s_Energy_Bin_Pos_102;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_102 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_102;   
  
  Energy_Bin_Pos_103 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_103   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_103 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E103_C1_L_Pos and PEAK_C1_Pos <= s_E103_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_103 <= s_Energy_Bin_Pos_103 +'1';
		 Energy_Bin_Pos_Rdy_103 <= '1';
		else
		 s_Energy_Bin_Pos_103 <= s_Energy_Bin_Pos_103;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_103 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_103;   
  
  Energy_Bin_Pos_104 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_104   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_104 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E104_C1_L_Pos and PEAK_C1_Pos <= s_E104_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_104 <= s_Energy_Bin_Pos_104 +'1';
		 Energy_Bin_Pos_Rdy_104 <= '1';
		else
		 s_Energy_Bin_Pos_104 <= s_Energy_Bin_Pos_104;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_104 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_104;   
 
 
  Energy_Bin_Pos_105 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_105   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_105 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E105_C1_L_Pos and PEAK_C1_Pos <= s_E105_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_105 <= s_Energy_Bin_Pos_105 +'1';
		 Energy_Bin_Pos_Rdy_105 <= '1';
		else
		 s_Energy_Bin_Pos_105 <= s_Energy_Bin_Pos_105;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_105 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_105;  
 
  
  Energy_Bin_Pos_106 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_106   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_106 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E106_C1_L_Pos and PEAK_C1_Pos <= s_E106_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_106 <= s_Energy_Bin_Pos_106 +'1';
		 Energy_Bin_Pos_Rdy_106 <= '1';
		else
		 s_Energy_Bin_Pos_106 <= s_Energy_Bin_Pos_106;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_106 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_106;   
  
 Energy_Bin_Pos_107 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_107   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_107 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E107_C1_L_Pos and PEAK_C1_Pos <= s_E107_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_107 <= s_Energy_Bin_Pos_107 +'1';
		 Energy_Bin_Pos_Rdy_107 <= '1';
		else
		 s_Energy_Bin_Pos_107 <= s_Energy_Bin_Pos_107;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_107 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_107;   
  
  Energy_Bin_Pos_108 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_108   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_108 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E108_C1_L_Pos and PEAK_C1_Pos <= s_E108_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_108 <= s_Energy_Bin_Pos_108 +'1';
		 Energy_Bin_Pos_Rdy_108 <= '1';
		else
		 s_Energy_Bin_Pos_108 <= s_Energy_Bin_Pos_108;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_108 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_108;   
  
  Energy_Bin_Pos_109 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_109   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_109 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E109_C1_L_Pos and PEAK_C1_Pos <= s_E109_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_109 <= s_Energy_Bin_Pos_109 +'1';
		 Energy_Bin_Pos_Rdy_109 <= '1';
		else
		 s_Energy_Bin_Pos_109 <= s_Energy_Bin_Pos_109;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_109 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_109;     
  
     Energy_Bin_Pos_110 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_110   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_110 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E110_C1_L_Pos and PEAK_C1_Pos <= s_E110_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_110 <= s_Energy_Bin_Pos_110 +'1';
		 Energy_Bin_Pos_Rdy_110 <= '1';
		else
		 s_Energy_Bin_Pos_110 <= s_Energy_Bin_Pos_110;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_110 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_110;    
  
  Energy_Bin_Pos_111 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_111   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_111 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E111_C1_L_Pos and PEAK_C1_Pos <= s_E111_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_111 <= s_Energy_Bin_Pos_111 +'1';
		 Energy_Bin_Pos_Rdy_111 <= '1';
		else
		 s_Energy_Bin_Pos_111 <= s_Energy_Bin_Pos_111;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_111 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_111;   
  
  Energy_Bin_Pos_112 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_112   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_112 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E112_C1_L_Pos and PEAK_C1_Pos <= s_E112_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_112 <= s_Energy_Bin_Pos_112 +'1';
		 Energy_Bin_Pos_Rdy_112 <= '1';
		else
		 s_Energy_Bin_Pos_112 <= s_Energy_Bin_Pos_112;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_112 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_112;   
  
  Energy_Bin_Pos_113 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_113   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_113 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E113_C1_L_Pos and PEAK_C1_Pos <= s_E113_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_113 <= s_Energy_Bin_Pos_113 +'1';
		 Energy_Bin_Pos_Rdy_113 <= '1';
		else
		 s_Energy_Bin_Pos_113 <= s_Energy_Bin_Pos_113;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_113 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_113;   
  
  Energy_Bin_Pos_114 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_114   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_114 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E114_C1_L_Pos and PEAK_C1_Pos <= s_E114_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_114 <= s_Energy_Bin_Pos_114 +'1';
		 Energy_Bin_Pos_Rdy_114 <= '1';
		else
		 s_Energy_Bin_Pos_114 <= s_Energy_Bin_Pos_114;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_114 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_114;   
 
 
  Energy_Bin_Pos_115 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_115   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_115 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E115_C1_L_Pos and PEAK_C1_Pos <= s_E115_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_115 <= s_Energy_Bin_Pos_115 +'1';
		 Energy_Bin_Pos_Rdy_115 <= '1';
		else
		 s_Energy_Bin_Pos_115 <= s_Energy_Bin_Pos_115;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_115 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_115;  
 
  
  Energy_Bin_Pos_116 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_116   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_116 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E116_C1_L_Pos and PEAK_C1_Pos <= s_E116_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_116 <= s_Energy_Bin_Pos_116 +'1';
		 Energy_Bin_Pos_Rdy_116 <= '1';
		else
		 s_Energy_Bin_Pos_116 <= s_Energy_Bin_Pos_116;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_116 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_116;   
  
 Energy_Bin_Pos_117 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_117   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_117 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E117_C1_L_Pos and PEAK_C1_Pos <= s_E117_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_117 <= s_Energy_Bin_Pos_117 +'1';
		 Energy_Bin_Pos_Rdy_117 <= '1';
		else
		 s_Energy_Bin_Pos_117 <= s_Energy_Bin_Pos_117;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_117 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_117;   
  
  Energy_Bin_Pos_118 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_118   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_118 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E118_C1_L_Pos and PEAK_C1_Pos <= s_E118_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_118 <= s_Energy_Bin_Pos_118 +'1';
		 Energy_Bin_Pos_Rdy_118 <= '1';
		else
		 s_Energy_Bin_Pos_118 <= s_Energy_Bin_Pos_118;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_118 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_118;   
  
  Energy_Bin_Pos_119 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_119   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_119 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E119_C1_L_Pos and PEAK_C1_Pos <= s_E119_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_119 <= s_Energy_Bin_Pos_119 +'1';
		 Energy_Bin_Pos_Rdy_119 <= '1';
		else
		 s_Energy_Bin_Pos_119 <= s_Energy_Bin_Pos_119;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_119 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_119;      
  
     Energy_Bin_Pos_120 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_120   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_120 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E120_C1_L_Pos and PEAK_C1_Pos <= s_E120_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_120 <= s_Energy_Bin_Pos_120 +'1';
		 Energy_Bin_Pos_Rdy_120 <= '1';
		else
		 s_Energy_Bin_Pos_120 <= s_Energy_Bin_Pos_120;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_120 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_120;    
  
  Energy_Bin_Pos_121 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_121   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_121 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E121_C1_L_Pos and PEAK_C1_Pos <= s_E121_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_121 <= s_Energy_Bin_Pos_121 +'1';
		 Energy_Bin_Pos_Rdy_121 <= '1';
		else
		 s_Energy_Bin_Pos_121 <= s_Energy_Bin_Pos_121;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_121 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_121;   
  
  Energy_Bin_Pos_122 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_122   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_122 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E122_C1_L_Pos and PEAK_C1_Pos <= s_E122_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_122 <= s_Energy_Bin_Pos_122 +'1';
		 Energy_Bin_Pos_Rdy_122 <= '1';
		else
		 s_Energy_Bin_Pos_122 <= s_Energy_Bin_Pos_122;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_122 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_122;   
  
  Energy_Bin_Pos_123 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_123   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_123 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E123_C1_L_Pos and PEAK_C1_Pos <= s_E123_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_123 <= s_Energy_Bin_Pos_123 +'1';
		 Energy_Bin_Pos_Rdy_123 <= '1';
		else
		 s_Energy_Bin_Pos_123 <= s_Energy_Bin_Pos_123;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_123 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_123;   
  
  Energy_Bin_Pos_124 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_124   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_124 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E124_C1_L_Pos and PEAK_C1_Pos <= s_E124_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_124 <= s_Energy_Bin_Pos_124 +'1';
		 Energy_Bin_Pos_Rdy_124 <= '1';
		else
		 s_Energy_Bin_Pos_124 <= s_Energy_Bin_Pos_124;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_124 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_124;   
 
 
  Energy_Bin_Pos_125 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_125   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_125 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E125_C1_L_Pos and PEAK_C1_Pos <= s_E125_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_125 <= s_Energy_Bin_Pos_125 +'1';
		 Energy_Bin_Pos_Rdy_125 <= '1';
		else
		 s_Energy_Bin_Pos_125 <= s_Energy_Bin_Pos_125;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_125 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_125;  
 
  
  Energy_Bin_Pos_126 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_126   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_126 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E126_C1_L_Pos and PEAK_C1_Pos <= s_E126_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_126 <= s_Energy_Bin_Pos_126 +'1';
		 Energy_Bin_Pos_Rdy_126 <= '1';
		else
		 s_Energy_Bin_Pos_126 <= s_Energy_Bin_Pos_126;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_126 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_126;   
  
 Energy_Bin_Pos_127 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_127   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_127 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E127_C1_L_Pos and PEAK_C1_Pos <= s_E127_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_127 <= s_Energy_Bin_Pos_127 +'1';
		 Energy_Bin_Pos_Rdy_127 <= '1';
		else
		 s_Energy_Bin_Pos_127 <= s_Energy_Bin_Pos_127;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_127 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_127;   
  
  Energy_Bin_Pos_128 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_128   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_128 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E128_C1_L_Pos and PEAK_C1_Pos <= s_E128_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_128 <= s_Energy_Bin_Pos_128 +'1';
		 Energy_Bin_Pos_Rdy_128 <= '1';
		else
		 s_Energy_Bin_Pos_128 <= s_Energy_Bin_Pos_128;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_128 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_128;   
  
  Energy_Bin_Pos_129 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_129   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_129 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E129_C1_L_Pos and PEAK_C1_Pos <= s_E129_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_129 <= s_Energy_Bin_Pos_129 +'1';
		 Energy_Bin_Pos_Rdy_129 <= '1';
		else
		 s_Energy_Bin_Pos_129 <= s_Energy_Bin_Pos_129;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_129 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_129;       
  
     Energy_Bin_Pos_130 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_130   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_130 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E130_C1_L_Pos and PEAK_C1_Pos <= s_E130_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_130 <= s_Energy_Bin_Pos_130 +'1';
		 Energy_Bin_Pos_Rdy_130 <= '1';
		else
		 s_Energy_Bin_Pos_130 <= s_Energy_Bin_Pos_130;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_130 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_130;    
  
  Energy_Bin_Pos_131 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_131   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_131 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E131_C1_L_Pos and PEAK_C1_Pos <= s_E131_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_131 <= s_Energy_Bin_Pos_131 +'1';
		 Energy_Bin_Pos_Rdy_131 <= '1';
		else
		 s_Energy_Bin_Pos_131 <= s_Energy_Bin_Pos_131;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_131 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_131;   
  
  Energy_Bin_Pos_132 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_132   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_132 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E132_C1_L_Pos and PEAK_C1_Pos <= s_E132_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_132 <= s_Energy_Bin_Pos_132 +'1';
		 Energy_Bin_Pos_Rdy_132 <= '1';
		else
		 s_Energy_Bin_Pos_132 <= s_Energy_Bin_Pos_132;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_132 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_132;   
  
  Energy_Bin_Pos_133 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_133   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_133 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E133_C1_L_Pos and PEAK_C1_Pos <= s_E133_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_133 <= s_Energy_Bin_Pos_133 +'1';
		 Energy_Bin_Pos_Rdy_133 <= '1';
		else
		 s_Energy_Bin_Pos_133 <= s_Energy_Bin_Pos_133;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_133 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_133;   
  
  Energy_Bin_Pos_134 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_134   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_134 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E134_C1_L_Pos and PEAK_C1_Pos <= s_E134_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_134 <= s_Energy_Bin_Pos_134 +'1';
		 Energy_Bin_Pos_Rdy_134 <= '1';
		else
		 s_Energy_Bin_Pos_134 <= s_Energy_Bin_Pos_134;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_134 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_134;   
 
 
  Energy_Bin_Pos_135 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_135   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_135 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E135_C1_L_Pos and PEAK_C1_Pos <= s_E135_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_135 <= s_Energy_Bin_Pos_135 +'1';
		 Energy_Bin_Pos_Rdy_135 <= '1';
		else
		 s_Energy_Bin_Pos_135 <= s_Energy_Bin_Pos_135;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_135 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_135;  
 
  
  Energy_Bin_Pos_136 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_136   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_136 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E136_C1_L_Pos and PEAK_C1_Pos <= s_E136_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_136 <= s_Energy_Bin_Pos_136 +'1';
		 Energy_Bin_Pos_Rdy_136 <= '1';
		else
		 s_Energy_Bin_Pos_136 <= s_Energy_Bin_Pos_136;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_136 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_136;   
  
 Energy_Bin_Pos_137 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_137   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_137 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E137_C1_L_Pos and PEAK_C1_Pos <= s_E137_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_137 <= s_Energy_Bin_Pos_137 +'1';
		 Energy_Bin_Pos_Rdy_137 <= '1';
		else
		 s_Energy_Bin_Pos_137 <= s_Energy_Bin_Pos_137;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_137 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_137;   
  
  Energy_Bin_Pos_138 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_138   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_138 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E138_C1_L_Pos and PEAK_C1_Pos <= s_E138_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_138 <= s_Energy_Bin_Pos_138 +'1';
		 Energy_Bin_Pos_Rdy_138 <= '1';
		else
		 s_Energy_Bin_Pos_138 <= s_Energy_Bin_Pos_138;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_138 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_138;   
  
  Energy_Bin_Pos_139 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_139   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_139 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E139_C1_L_Pos and PEAK_C1_Pos <= s_E139_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_139 <= s_Energy_Bin_Pos_139 +'1';
		 Energy_Bin_Pos_Rdy_139 <= '1';
		else
		 s_Energy_Bin_Pos_139 <= s_Energy_Bin_Pos_139;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_139 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_139;         
  
     Energy_Bin_Pos_140 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_140   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_140 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E140_C1_L_Pos and PEAK_C1_Pos <= s_E140_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_140 <= s_Energy_Bin_Pos_140 +'1';
		 Energy_Bin_Pos_Rdy_140 <= '1';
		else
		 s_Energy_Bin_Pos_140 <= s_Energy_Bin_Pos_140;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_140 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_140;    
  
  Energy_Bin_Pos_141 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_141   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_141 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E141_C1_L_Pos and PEAK_C1_Pos <= s_E141_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_141 <= s_Energy_Bin_Pos_141 +'1';
		 Energy_Bin_Pos_Rdy_141 <= '1';
		else
		 s_Energy_Bin_Pos_141 <= s_Energy_Bin_Pos_141;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_141 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_141;   
  
  Energy_Bin_Pos_142 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_142   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_142 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E142_C1_L_Pos and PEAK_C1_Pos <= s_E142_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_142 <= s_Energy_Bin_Pos_142 +'1';
		 Energy_Bin_Pos_Rdy_142 <= '1';
		else
		 s_Energy_Bin_Pos_142 <= s_Energy_Bin_Pos_142;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_142 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_142;   
  
  Energy_Bin_Pos_143 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_143   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_143 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E143_C1_L_Pos and PEAK_C1_Pos <= s_E143_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_143 <= s_Energy_Bin_Pos_143 +'1';
		 Energy_Bin_Pos_Rdy_143 <= '1';
		else
		 s_Energy_Bin_Pos_143 <= s_Energy_Bin_Pos_143;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_143 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_143;   
  
  Energy_Bin_Pos_144 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_144   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_144 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E144_C1_L_Pos and PEAK_C1_Pos <= s_E144_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_144 <= s_Energy_Bin_Pos_144 +'1';
		 Energy_Bin_Pos_Rdy_144 <= '1';
		else
		 s_Energy_Bin_Pos_144 <= s_Energy_Bin_Pos_144;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_144 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_144;   
 
 
  Energy_Bin_Pos_145 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_145   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_145 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E145_C1_L_Pos and PEAK_C1_Pos <= s_E145_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_145 <= s_Energy_Bin_Pos_145 +'1';
		 Energy_Bin_Pos_Rdy_145 <= '1';
		else
		 s_Energy_Bin_Pos_145 <= s_Energy_Bin_Pos_145;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_145 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_145;  
 
  
  Energy_Bin_Pos_146 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_146   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_146 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E146_C1_L_Pos and PEAK_C1_Pos <= s_E146_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_146 <= s_Energy_Bin_Pos_146 +'1';
		 Energy_Bin_Pos_Rdy_146 <= '1';
		else
		 s_Energy_Bin_Pos_146 <= s_Energy_Bin_Pos_146;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_146 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_146;   
  
 Energy_Bin_Pos_147 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_147   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_147 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E147_C1_L_Pos and PEAK_C1_Pos <= s_E147_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_147 <= s_Energy_Bin_Pos_147 +'1';
		 Energy_Bin_Pos_Rdy_147 <= '1';
		else
		 s_Energy_Bin_Pos_147 <= s_Energy_Bin_Pos_147;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_147 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_147;   
  
  Energy_Bin_Pos_148 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_148   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_148 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E148_C1_L_Pos and PEAK_C1_Pos <= s_E148_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_148 <= s_Energy_Bin_Pos_148 +'1';
		 Energy_Bin_Pos_Rdy_148 <= '1';
		else
		 s_Energy_Bin_Pos_148 <= s_Energy_Bin_Pos_148;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_148 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_148;   
  
  Energy_Bin_Pos_149 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_149   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_149 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E149_C1_L_Pos and PEAK_C1_Pos <= s_E149_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_149 <= s_Energy_Bin_Pos_149 +'1';
		 Energy_Bin_Pos_Rdy_149 <= '1';
		else
		 s_Energy_Bin_Pos_149 <= s_Energy_Bin_Pos_149;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_149 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_149;          
  
  
     Energy_Bin_Pos_150 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_150   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_150 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E150_C1_L_Pos and PEAK_C1_Pos <= s_E150_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_150 <= s_Energy_Bin_Pos_150 +'1';
		 Energy_Bin_Pos_Rdy_150 <= '1';
		else
		 s_Energy_Bin_Pos_150 <= s_Energy_Bin_Pos_150;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_150 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_150;    
  
  Energy_Bin_Pos_151 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_151   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_151 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E151_C1_L_Pos and PEAK_C1_Pos <= s_E151_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_151 <= s_Energy_Bin_Pos_151 +'1';
		 Energy_Bin_Pos_Rdy_151 <= '1';
		else
		 s_Energy_Bin_Pos_151 <= s_Energy_Bin_Pos_151;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_151 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_151;   
  
  Energy_Bin_Pos_152 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_152   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_152 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E152_C1_L_Pos and PEAK_C1_Pos <= s_E152_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_152 <= s_Energy_Bin_Pos_152 +'1';
		 Energy_Bin_Pos_Rdy_152 <= '1';
		else
		 s_Energy_Bin_Pos_152 <= s_Energy_Bin_Pos_152;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_152 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_152;   
  
  Energy_Bin_Pos_153 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_153   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_153 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E153_C1_L_Pos and PEAK_C1_Pos <= s_E153_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_153 <= s_Energy_Bin_Pos_153 +'1';
		 Energy_Bin_Pos_Rdy_153 <= '1';
		else
		 s_Energy_Bin_Pos_153 <= s_Energy_Bin_Pos_153;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_153 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_153;   
  
  Energy_Bin_Pos_154 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_154   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_154 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E154_C1_L_Pos and PEAK_C1_Pos <= s_E154_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_154 <= s_Energy_Bin_Pos_154 +'1';
		 Energy_Bin_Pos_Rdy_154 <= '1';
		else
		 s_Energy_Bin_Pos_154 <= s_Energy_Bin_Pos_154;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_154 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_154;   
 
 
  Energy_Bin_Pos_155 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_155   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_155 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E155_C1_L_Pos and PEAK_C1_Pos <= s_E155_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_155 <= s_Energy_Bin_Pos_155 +'1';
		 Energy_Bin_Pos_Rdy_155 <= '1';
		else
		 s_Energy_Bin_Pos_155 <= s_Energy_Bin_Pos_155;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_155 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_155;  
 
  
  Energy_Bin_Pos_156 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_156   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_156 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E156_C1_L_Pos and PEAK_C1_Pos <= s_E156_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_156 <= s_Energy_Bin_Pos_156 +'1';
		 Energy_Bin_Pos_Rdy_156 <= '1';
		else
		 s_Energy_Bin_Pos_156 <= s_Energy_Bin_Pos_156;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_156 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_156;   
  
 Energy_Bin_Pos_157 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_157   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_157 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E157_C1_L_Pos and PEAK_C1_Pos <= s_E157_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_157 <= s_Energy_Bin_Pos_157 +'1';
		 Energy_Bin_Pos_Rdy_157 <= '1';
		else
		 s_Energy_Bin_Pos_157 <= s_Energy_Bin_Pos_157;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_157 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_157;   
  
  Energy_Bin_Pos_158 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_158   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_158 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E158_C1_L_Pos and PEAK_C1_Pos <= s_E158_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_158 <= s_Energy_Bin_Pos_158 +'1';
		 Energy_Bin_Pos_Rdy_158 <= '1';
		else
		 s_Energy_Bin_Pos_158 <= s_Energy_Bin_Pos_158;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_158 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_158;   
  
  Energy_Bin_Pos_159 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_159   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_159 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E159_C1_L_Pos and PEAK_C1_Pos <= s_E159_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_159 <= s_Energy_Bin_Pos_159 +'1';
		 Energy_Bin_Pos_Rdy_159 <= '1';
		else
		 s_Energy_Bin_Pos_159 <= s_Energy_Bin_Pos_159;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_159 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_159;           
  
     Energy_Bin_Pos_160 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_160   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_160 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E160_C1_L_Pos and PEAK_C1_Pos <= s_E160_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_160 <= s_Energy_Bin_Pos_160 +'1';
		 Energy_Bin_Pos_Rdy_160 <= '1';
		else
		 s_Energy_Bin_Pos_160 <= s_Energy_Bin_Pos_160;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_160 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_160;    
  
  Energy_Bin_Pos_161 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_161   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_161 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E161_C1_L_Pos and PEAK_C1_Pos <= s_E161_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_161 <= s_Energy_Bin_Pos_161 +'1';
		 Energy_Bin_Pos_Rdy_161 <= '1';
		else
		 s_Energy_Bin_Pos_161 <= s_Energy_Bin_Pos_161;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_161 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_161;   
  
  Energy_Bin_Pos_162 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_162   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_162 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E162_C1_L_Pos and PEAK_C1_Pos <= s_E162_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_162 <= s_Energy_Bin_Pos_162 +'1';
		 Energy_Bin_Pos_Rdy_162 <= '1';
		else
		 s_Energy_Bin_Pos_162 <= s_Energy_Bin_Pos_162;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_162 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_162;   
  
  Energy_Bin_Pos_163 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_163   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_163 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E163_C1_L_Pos and PEAK_C1_Pos <= s_E163_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_163 <= s_Energy_Bin_Pos_163 +'1';
		 Energy_Bin_Pos_Rdy_163 <= '1';
		else
		 s_Energy_Bin_Pos_163 <= s_Energy_Bin_Pos_163;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_163 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_163;   
  
  Energy_Bin_Pos_164 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_164   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_164 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E164_C1_L_Pos and PEAK_C1_Pos <= s_E164_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_164 <= s_Energy_Bin_Pos_164 +'1';
		 Energy_Bin_Pos_Rdy_164 <= '1';
		else
		 s_Energy_Bin_Pos_164 <= s_Energy_Bin_Pos_164;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_164 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_164;   
 
 
  Energy_Bin_Pos_165 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_165   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_165 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E165_C1_L_Pos and PEAK_C1_Pos <= s_E165_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_165 <= s_Energy_Bin_Pos_165 +'1';
		 Energy_Bin_Pos_Rdy_165 <= '1';
		else
		 s_Energy_Bin_Pos_165 <= s_Energy_Bin_Pos_165;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_165 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_165;  
 
  
  Energy_Bin_Pos_166 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_166   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_166 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E166_C1_L_Pos and PEAK_C1_Pos <= s_E166_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_166 <= s_Energy_Bin_Pos_166 +'1';
		 Energy_Bin_Pos_Rdy_166 <= '1';
		else
		 s_Energy_Bin_Pos_166 <= s_Energy_Bin_Pos_166;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_166 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_166;   
  
 Energy_Bin_Pos_167 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_167   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_167 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E167_C1_L_Pos and PEAK_C1_Pos <= s_E167_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_167 <= s_Energy_Bin_Pos_167 +'1';
		 Energy_Bin_Pos_Rdy_167 <= '1';
		else
		 s_Energy_Bin_Pos_167 <= s_Energy_Bin_Pos_167;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_167 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_167;   
  
  Energy_Bin_Pos_168 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_168   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_168 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E168_C1_L_Pos and PEAK_C1_Pos <= s_E168_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_168 <= s_Energy_Bin_Pos_168 +'1';
		 Energy_Bin_Pos_Rdy_168 <= '1';
		else
		 s_Energy_Bin_Pos_168 <= s_Energy_Bin_Pos_168;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_168 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_168;   
  
  Energy_Bin_Pos_169 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_169   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_169 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E169_C1_L_Pos and PEAK_C1_Pos <= s_E169_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_169 <= s_Energy_Bin_Pos_169 +'1';
		 Energy_Bin_Pos_Rdy_169 <= '1';
		else
		 s_Energy_Bin_Pos_169 <= s_Energy_Bin_Pos_169;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_169 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_169;         
  
     Energy_Bin_Pos_170 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_170   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_170 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E170_C1_L_Pos and PEAK_C1_Pos <= s_E170_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_170 <= s_Energy_Bin_Pos_170 +'1';
		 Energy_Bin_Pos_Rdy_170 <= '1';
		else
		 s_Energy_Bin_Pos_170 <= s_Energy_Bin_Pos_170;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_170 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_170;    
  
  Energy_Bin_Pos_171 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_171   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_171 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E171_C1_L_Pos and PEAK_C1_Pos <= s_E171_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_171 <= s_Energy_Bin_Pos_171 +'1';
		 Energy_Bin_Pos_Rdy_171 <= '1';
		else
		 s_Energy_Bin_Pos_171 <= s_Energy_Bin_Pos_171;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_171 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_171;   
  
  Energy_Bin_Pos_172 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_172   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_172 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E172_C1_L_Pos and PEAK_C1_Pos <= s_E172_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_172 <= s_Energy_Bin_Pos_172 +'1';
		 Energy_Bin_Pos_Rdy_172 <= '1';
		else
		 s_Energy_Bin_Pos_172 <= s_Energy_Bin_Pos_172;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_172 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_172;   
  
  Energy_Bin_Pos_173 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_173   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_173 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E173_C1_L_Pos and PEAK_C1_Pos <= s_E173_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_173 <= s_Energy_Bin_Pos_173 +'1';
		 Energy_Bin_Pos_Rdy_173 <= '1';
		else
		 s_Energy_Bin_Pos_173 <= s_Energy_Bin_Pos_173;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_173 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_173;   
  
  Energy_Bin_Pos_174 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_174   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_174 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E174_C1_L_Pos and PEAK_C1_Pos <= s_E174_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_174 <= s_Energy_Bin_Pos_174 +'1';
		 Energy_Bin_Pos_Rdy_174 <= '1';
		else
		 s_Energy_Bin_Pos_174 <= s_Energy_Bin_Pos_174;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_174 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_174;   
 
 
  Energy_Bin_Pos_175 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_175   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_175 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E175_C1_L_Pos and PEAK_C1_Pos <= s_E175_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_175 <= s_Energy_Bin_Pos_175 +'1';
		 Energy_Bin_Pos_Rdy_175 <= '1';
		else
		 s_Energy_Bin_Pos_175 <= s_Energy_Bin_Pos_175;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_175 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_175;  
 
  
  Energy_Bin_Pos_176 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_176   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_176 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E176_C1_L_Pos and PEAK_C1_Pos <= s_E176_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_176 <= s_Energy_Bin_Pos_176 +'1';
		 Energy_Bin_Pos_Rdy_176 <= '1';
		else
		 s_Energy_Bin_Pos_176 <= s_Energy_Bin_Pos_176;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_176 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_176;   
  
 Energy_Bin_Pos_177 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_177   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_177 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E177_C1_L_Pos and PEAK_C1_Pos <= s_E177_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_177 <= s_Energy_Bin_Pos_177 +'1';
		 Energy_Bin_Pos_Rdy_177 <= '1';
		else
		 s_Energy_Bin_Pos_177 <= s_Energy_Bin_Pos_177;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_177 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_177;   
  
  Energy_Bin_Pos_178 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_178   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_178 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E178_C1_L_Pos and PEAK_C1_Pos <= s_E178_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_178 <= s_Energy_Bin_Pos_178 +'1';
		 Energy_Bin_Pos_Rdy_178 <= '1';
		else
		 s_Energy_Bin_Pos_178 <= s_Energy_Bin_Pos_178;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_178 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_178;   
  
  Energy_Bin_Pos_179 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_179   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_179 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E179_C1_L_Pos and PEAK_C1_Pos <= s_E179_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_179 <= s_Energy_Bin_Pos_179 +'1';
		 Energy_Bin_Pos_Rdy_179 <= '1';
		else
		 s_Energy_Bin_Pos_179 <= s_Energy_Bin_Pos_179;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_179 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_179;       
  
     Energy_Bin_Pos_180 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_180   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_180 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E180_C1_L_Pos and PEAK_C1_Pos <= s_E180_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_180 <= s_Energy_Bin_Pos_180 +'1';
		 Energy_Bin_Pos_Rdy_180 <= '1';
		else
		 s_Energy_Bin_Pos_180 <= s_Energy_Bin_Pos_180;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_180 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_180;    
  
  Energy_Bin_Pos_181 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_181   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_181 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E181_C1_L_Pos and PEAK_C1_Pos <= s_E181_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_181 <= s_Energy_Bin_Pos_181 +'1';
		 Energy_Bin_Pos_Rdy_181 <= '1';
		else
		 s_Energy_Bin_Pos_181 <= s_Energy_Bin_Pos_181;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_181 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_181;   
  
  Energy_Bin_Pos_182 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_182   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_182 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E182_C1_L_Pos and PEAK_C1_Pos <= s_E182_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_182 <= s_Energy_Bin_Pos_182 +'1';
		 Energy_Bin_Pos_Rdy_182 <= '1';
		else
		 s_Energy_Bin_Pos_182 <= s_Energy_Bin_Pos_182;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_182 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_182;   
  
  Energy_Bin_Pos_183 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_183   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_183 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E183_C1_L_Pos and PEAK_C1_Pos <= s_E183_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_183 <= s_Energy_Bin_Pos_183 +'1';
		 Energy_Bin_Pos_Rdy_183 <= '1';
		else
		 s_Energy_Bin_Pos_183 <= s_Energy_Bin_Pos_183;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_183 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_183;   
  
  Energy_Bin_Pos_184 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_184   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_184 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E184_C1_L_Pos and PEAK_C1_Pos <= s_E184_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_184 <= s_Energy_Bin_Pos_184 +'1';
		 Energy_Bin_Pos_Rdy_184 <= '1';
		else
		 s_Energy_Bin_Pos_184 <= s_Energy_Bin_Pos_184;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_184 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_184;   
 
 
  Energy_Bin_Pos_185 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_185   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_185 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E185_C1_L_Pos and PEAK_C1_Pos <= s_E185_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_185 <= s_Energy_Bin_Pos_185 +'1';
		 Energy_Bin_Pos_Rdy_185 <= '1';
		else
		 s_Energy_Bin_Pos_185 <= s_Energy_Bin_Pos_185;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_185 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_185;  
 
  
  Energy_Bin_Pos_186 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_186   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_186 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E186_C1_L_Pos and PEAK_C1_Pos <= s_E186_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_186 <= s_Energy_Bin_Pos_186 +'1';
		 Energy_Bin_Pos_Rdy_186 <= '1';
		else
		 s_Energy_Bin_Pos_186 <= s_Energy_Bin_Pos_186;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_186 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_186;   
  
 Energy_Bin_Pos_187 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_187   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_187 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E187_C1_L_Pos and PEAK_C1_Pos <= s_E187_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_187 <= s_Energy_Bin_Pos_187 +'1';
		 Energy_Bin_Pos_Rdy_187 <= '1';
		else
		 s_Energy_Bin_Pos_187 <= s_Energy_Bin_Pos_187;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_187 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_187;   
  
  Energy_Bin_Pos_188 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_188   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_188 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E188_C1_L_Pos and PEAK_C1_Pos <= s_E188_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_188 <= s_Energy_Bin_Pos_188 +'1';
		 Energy_Bin_Pos_Rdy_188 <= '1';
		else
		 s_Energy_Bin_Pos_188 <= s_Energy_Bin_Pos_188;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_188 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_188;   
  
  Energy_Bin_Pos_189 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_189   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_189 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E189_C1_L_Pos and PEAK_C1_Pos <= s_E189_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_189 <= s_Energy_Bin_Pos_189 +'1';
		 Energy_Bin_Pos_Rdy_189 <= '1';
		else
		 s_Energy_Bin_Pos_189 <= s_Energy_Bin_Pos_189;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_189 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_189;      
  
     Energy_Bin_Pos_190 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_190   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_190 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E190_C1_L_Pos and PEAK_C1_Pos <= s_E190_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_190 <= s_Energy_Bin_Pos_190 +'1';
		 Energy_Bin_Pos_Rdy_190 <= '1';
		else
		 s_Energy_Bin_Pos_190 <= s_Energy_Bin_Pos_190;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_190 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_190;    
  
  Energy_Bin_Pos_191 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_191   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_191 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E191_C1_L_Pos and PEAK_C1_Pos <= s_E191_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_191 <= s_Energy_Bin_Pos_191 +'1';
		 Energy_Bin_Pos_Rdy_191 <= '1';
		else
		 s_Energy_Bin_Pos_191 <= s_Energy_Bin_Pos_191;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_191 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_191;   
  
  Energy_Bin_Pos_192 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_192   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_192 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E192_C1_L_Pos and PEAK_C1_Pos <= s_E192_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_192 <= s_Energy_Bin_Pos_192 +'1';
		 Energy_Bin_Pos_Rdy_192 <= '1';
		else
		 s_Energy_Bin_Pos_192 <= s_Energy_Bin_Pos_192;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_192 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_192;   
  
  Energy_Bin_Pos_193 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_193   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_193 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E193_C1_L_Pos and PEAK_C1_Pos <= s_E193_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_193 <= s_Energy_Bin_Pos_193 +'1';
		 Energy_Bin_Pos_Rdy_193 <= '1';
		else
		 s_Energy_Bin_Pos_193 <= s_Energy_Bin_Pos_193;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_193 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_193;   
  
  Energy_Bin_Pos_194 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_194   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_194 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E194_C1_L_Pos and PEAK_C1_Pos <= s_E194_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_194 <= s_Energy_Bin_Pos_194 +'1';
		 Energy_Bin_Pos_Rdy_194 <= '1';
		else
		 s_Energy_Bin_Pos_194 <= s_Energy_Bin_Pos_194;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_194 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_194;   
 
 
  Energy_Bin_Pos_195 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_195   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_195 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E195_C1_L_Pos and PEAK_C1_Pos <= s_E195_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_195 <= s_Energy_Bin_Pos_195 +'1';
		 Energy_Bin_Pos_Rdy_195 <= '1';
		else
		 s_Energy_Bin_Pos_195 <= s_Energy_Bin_Pos_195;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_195 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_195;  
 
  
  Energy_Bin_Pos_196 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_196   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_196 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E196_C1_L_Pos and PEAK_C1_Pos <= s_E196_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_196 <= s_Energy_Bin_Pos_196 +'1';
		 Energy_Bin_Pos_Rdy_196 <= '1';
		else
		 s_Energy_Bin_Pos_196 <= s_Energy_Bin_Pos_196;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_196 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_196;   
  
 Energy_Bin_Pos_197 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_197   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_197 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E197_C1_L_Pos and PEAK_C1_Pos <= s_E197_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_197 <= s_Energy_Bin_Pos_197 +'1';
		 Energy_Bin_Pos_Rdy_197 <= '1';
		else
		 s_Energy_Bin_Pos_197 <= s_Energy_Bin_Pos_197;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_197 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_197;   
  
  Energy_Bin_Pos_198 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_198   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_198 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E198_C1_L_Pos and PEAK_C1_Pos <= s_E198_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_198 <= s_Energy_Bin_Pos_198 +'1';
		 Energy_Bin_Pos_Rdy_198 <= '1';
		else
		 s_Energy_Bin_Pos_198 <= s_Energy_Bin_Pos_198;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_198 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_198;   
  
  Energy_Bin_Pos_199 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_199   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_199 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E199_C1_L_Pos and PEAK_C1_Pos <= s_E199_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_199 <= s_Energy_Bin_Pos_199 +'1';
		 Energy_Bin_Pos_Rdy_199 <= '1';
		else
		 s_Energy_Bin_Pos_199 <= s_Energy_Bin_Pos_199;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_199 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_199;      
    
     Energy_Bin_Pos_200 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_200   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_200 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E200_C1_L_Pos and PEAK_C1_Pos <= s_E200_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_200 <= s_Energy_Bin_Pos_200 +'1';
		 Energy_Bin_Pos_Rdy_200 <= '1';
		else
		 s_Energy_Bin_Pos_200 <= s_Energy_Bin_Pos_200;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_200 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_200;    
  
  Energy_Bin_Pos_201 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_201   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_201 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E201_C1_L_Pos and PEAK_C1_Pos <= s_E201_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_201 <= s_Energy_Bin_Pos_201 +'1';
		 Energy_Bin_Pos_Rdy_201 <= '1';
		else
		 s_Energy_Bin_Pos_201 <= s_Energy_Bin_Pos_201;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_201 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_201;   
  
  Energy_Bin_Pos_202 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_202   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_202 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E202_C1_L_Pos and PEAK_C1_Pos <= s_E202_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_202 <= s_Energy_Bin_Pos_202 +'1';
		 Energy_Bin_Pos_Rdy_202 <= '1';
		else
		 s_Energy_Bin_Pos_202 <= s_Energy_Bin_Pos_202;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_202 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_202;   
  
  Energy_Bin_Pos_203 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_203   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_203 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E203_C1_L_Pos and PEAK_C1_Pos <= s_E203_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_203 <= s_Energy_Bin_Pos_203 +'1';
		 Energy_Bin_Pos_Rdy_203 <= '1';
		else
		 s_Energy_Bin_Pos_203 <= s_Energy_Bin_Pos_203;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_203 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_203;   
  
  Energy_Bin_Pos_204 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_204   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_204 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E204_C1_L_Pos and PEAK_C1_Pos <= s_E204_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_204 <= s_Energy_Bin_Pos_204 +'1';
		 Energy_Bin_Pos_Rdy_204 <= '1';
		else
		 s_Energy_Bin_Pos_204 <= s_Energy_Bin_Pos_204;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_204 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_204;   
 
 
  Energy_Bin_Pos_205 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_205   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_205 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E205_C1_L_Pos and PEAK_C1_Pos <= s_E205_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_205 <= s_Energy_Bin_Pos_205 +'1';
		 Energy_Bin_Pos_Rdy_205 <= '1';
		else
		 s_Energy_Bin_Pos_205 <= s_Energy_Bin_Pos_205;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_205 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_205;  
 
  
  Energy_Bin_Pos_206 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_206   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_206 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E206_C1_L_Pos and PEAK_C1_Pos <= s_E206_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_206 <= s_Energy_Bin_Pos_206 +'1';
		 Energy_Bin_Pos_Rdy_206 <= '1';
		else
		 s_Energy_Bin_Pos_206 <= s_Energy_Bin_Pos_206;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_206 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_206;   
  
 Energy_Bin_Pos_207 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_207   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_207 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E207_C1_L_Pos and PEAK_C1_Pos <= s_E207_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_207 <= s_Energy_Bin_Pos_207 +'1';
		 Energy_Bin_Pos_Rdy_207 <= '1';
		else
		 s_Energy_Bin_Pos_207 <= s_Energy_Bin_Pos_207;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_207 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_207;   
  
  Energy_Bin_Pos_208 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_208   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_208 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E208_C1_L_Pos and PEAK_C1_Pos <= s_E208_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_208 <= s_Energy_Bin_Pos_208 +'1';
		 Energy_Bin_Pos_Rdy_208 <= '1';
		else
		 s_Energy_Bin_Pos_208 <= s_Energy_Bin_Pos_208;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_208 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_208;   
  
  Energy_Bin_Pos_209 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_209   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_209 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E209_C1_L_Pos and PEAK_C1_Pos <= s_E209_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_209 <= s_Energy_Bin_Pos_209 +'1';
		 Energy_Bin_Pos_Rdy_209 <= '1';
		else
		 s_Energy_Bin_Pos_209 <= s_Energy_Bin_Pos_209;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_209 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_209;      
  
     Energy_Bin_Pos_210 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_210   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_210 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E210_C1_L_Pos and PEAK_C1_Pos <= s_E210_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_210 <= s_Energy_Bin_Pos_210 +'1';
		 Energy_Bin_Pos_Rdy_210 <= '1';
		else
		 s_Energy_Bin_Pos_210 <= s_Energy_Bin_Pos_210;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_210 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_210;    
  
  Energy_Bin_Pos_211 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_211   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_211 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E211_C1_L_Pos and PEAK_C1_Pos <= s_E211_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_211 <= s_Energy_Bin_Pos_211 +'1';
		 Energy_Bin_Pos_Rdy_211 <= '1';
		else
		 s_Energy_Bin_Pos_211 <= s_Energy_Bin_Pos_211;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_211 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_211;   
  
  Energy_Bin_Pos_212 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_212   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_212 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E212_C1_L_Pos and PEAK_C1_Pos <= s_E212_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_212 <= s_Energy_Bin_Pos_212 +'1';
		 Energy_Bin_Pos_Rdy_212 <= '1';
		else
		 s_Energy_Bin_Pos_212 <= s_Energy_Bin_Pos_212;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_212 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_212;   
  
  Energy_Bin_Pos_213 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_213   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_213 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E213_C1_L_Pos and PEAK_C1_Pos <= s_E213_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_213 <= s_Energy_Bin_Pos_213 +'1';
		 Energy_Bin_Pos_Rdy_213 <= '1';
		else
		 s_Energy_Bin_Pos_213 <= s_Energy_Bin_Pos_213;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_213 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_213;   
  
  Energy_Bin_Pos_214 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_214   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_214 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E214_C1_L_Pos and PEAK_C1_Pos <= s_E214_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_214 <= s_Energy_Bin_Pos_214 +'1';
		 Energy_Bin_Pos_Rdy_214 <= '1';
		else
		 s_Energy_Bin_Pos_214 <= s_Energy_Bin_Pos_214;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_214 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_214;   
 
 
  Energy_Bin_Pos_215 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_215   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_215 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E215_C1_L_Pos and PEAK_C1_Pos <= s_E215_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_215 <= s_Energy_Bin_Pos_215 +'1';
		 Energy_Bin_Pos_Rdy_215 <= '1';
		else
		 s_Energy_Bin_Pos_215 <= s_Energy_Bin_Pos_215;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_215 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_215;  
 
  
  Energy_Bin_Pos_216 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_216   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_216 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E216_C1_L_Pos and PEAK_C1_Pos <= s_E216_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_216 <= s_Energy_Bin_Pos_216 +'1';
		 Energy_Bin_Pos_Rdy_216 <= '1';
		else
		 s_Energy_Bin_Pos_216 <= s_Energy_Bin_Pos_216;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_216 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_216;   
  
 Energy_Bin_Pos_217 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_217   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_217 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E217_C1_L_Pos and PEAK_C1_Pos <= s_E217_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_217 <= s_Energy_Bin_Pos_217 +'1';
		 Energy_Bin_Pos_Rdy_217 <= '1';
		else
		 s_Energy_Bin_Pos_217 <= s_Energy_Bin_Pos_217;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_217 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_217;   
  
  Energy_Bin_Pos_218 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_218   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_218 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E218_C1_L_Pos and PEAK_C1_Pos <= s_E218_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_218 <= s_Energy_Bin_Pos_218 +'1';
		 Energy_Bin_Pos_Rdy_218 <= '1';
		else
		 s_Energy_Bin_Pos_218 <= s_Energy_Bin_Pos_218;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_218 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_218;   
  
  Energy_Bin_Pos_219 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_219   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_219 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E219_C1_L_Pos and PEAK_C1_Pos <= s_E219_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_219 <= s_Energy_Bin_Pos_219 +'1';
		 Energy_Bin_Pos_Rdy_219 <= '1';
		else
		 s_Energy_Bin_Pos_219 <= s_Energy_Bin_Pos_219;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_219 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_219;       
  
     Energy_Bin_Pos_220 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_220   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_220 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E220_C1_L_Pos and PEAK_C1_Pos <= s_E220_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_220 <= s_Energy_Bin_Pos_220 +'1';
		 Energy_Bin_Pos_Rdy_220 <= '1';
		else
		 s_Energy_Bin_Pos_220 <= s_Energy_Bin_Pos_220;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_220 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_220;    
  
  Energy_Bin_Pos_221 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_221   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_221 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E221_C1_L_Pos and PEAK_C1_Pos <= s_E221_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_221 <= s_Energy_Bin_Pos_221 +'1';
		 Energy_Bin_Pos_Rdy_221 <= '1';
		else
		 s_Energy_Bin_Pos_221 <= s_Energy_Bin_Pos_221;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_221 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_221;   
  
  Energy_Bin_Pos_222 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_222   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_222 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E222_C1_L_Pos and PEAK_C1_Pos <= s_E222_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_222 <= s_Energy_Bin_Pos_222 +'1';
		 Energy_Bin_Pos_Rdy_222 <= '1';
		else
		 s_Energy_Bin_Pos_222 <= s_Energy_Bin_Pos_222;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_222 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_222;   
  
  Energy_Bin_Pos_223 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_223   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_223 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E223_C1_L_Pos and PEAK_C1_Pos <= s_E223_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_223 <= s_Energy_Bin_Pos_223 +'1';
		 Energy_Bin_Pos_Rdy_223 <= '1';
		else
		 s_Energy_Bin_Pos_223 <= s_Energy_Bin_Pos_223;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_223 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_223;   
  
  Energy_Bin_Pos_224 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_224   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_224 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E224_C1_L_Pos and PEAK_C1_Pos <= s_E224_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_224 <= s_Energy_Bin_Pos_224 +'1';
		 Energy_Bin_Pos_Rdy_224 <= '1';
		else
		 s_Energy_Bin_Pos_224 <= s_Energy_Bin_Pos_224;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_224 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_224;   
 
 
  Energy_Bin_Pos_225 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_225   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_225 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E225_C1_L_Pos and PEAK_C1_Pos <= s_E225_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_225 <= s_Energy_Bin_Pos_225 +'1';
		 Energy_Bin_Pos_Rdy_225 <= '1';
		else
		 s_Energy_Bin_Pos_225 <= s_Energy_Bin_Pos_225;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_225 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_225;  
 
  
  Energy_Bin_Pos_226 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_226   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_226 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E226_C1_L_Pos and PEAK_C1_Pos <= s_E226_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_226 <= s_Energy_Bin_Pos_226 +'1';
		 Energy_Bin_Pos_Rdy_226 <= '1';
		else
		 s_Energy_Bin_Pos_226 <= s_Energy_Bin_Pos_226;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_226 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_226;   
  
 Energy_Bin_Pos_227 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_227   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_227 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E227_C1_L_Pos and PEAK_C1_Pos <= s_E227_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_227 <= s_Energy_Bin_Pos_227 +'1';
		 Energy_Bin_Pos_Rdy_227 <= '1';
		else
		 s_Energy_Bin_Pos_227 <= s_Energy_Bin_Pos_227;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_227 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_227;   
  
  Energy_Bin_Pos_228 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_228   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_228 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E228_C1_L_Pos and PEAK_C1_Pos <= s_E228_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_228 <= s_Energy_Bin_Pos_228 +'1';
		 Energy_Bin_Pos_Rdy_228 <= '1';
		else
		 s_Energy_Bin_Pos_228 <= s_Energy_Bin_Pos_228;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_228 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_228;   
  
  Energy_Bin_Pos_229 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_229   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_229 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E229_C1_L_Pos and PEAK_C1_Pos <= s_E229_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_229 <= s_Energy_Bin_Pos_229 +'1';
		 Energy_Bin_Pos_Rdy_229 <= '1';
		else
		 s_Energy_Bin_Pos_229 <= s_Energy_Bin_Pos_229;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_229 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_229;        
  
     Energy_Bin_Pos_230 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_230   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_230 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E230_C1_L_Pos and PEAK_C1_Pos <= s_E230_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_230 <= s_Energy_Bin_Pos_230 +'1';
		 Energy_Bin_Pos_Rdy_230 <= '1';
		else
		 s_Energy_Bin_Pos_230 <= s_Energy_Bin_Pos_230;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_230 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_230;    
  
  Energy_Bin_Pos_231 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_231   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_231 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E231_C1_L_Pos and PEAK_C1_Pos <= s_E231_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_231 <= s_Energy_Bin_Pos_231 +'1';
		 Energy_Bin_Pos_Rdy_231 <= '1';
		else
		 s_Energy_Bin_Pos_231 <= s_Energy_Bin_Pos_231;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_231 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_231;   
  
  Energy_Bin_Pos_232 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_232   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_232 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E232_C1_L_Pos and PEAK_C1_Pos <= s_E232_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_232 <= s_Energy_Bin_Pos_232 +'1';
		 Energy_Bin_Pos_Rdy_232 <= '1';
		else
		 s_Energy_Bin_Pos_232 <= s_Energy_Bin_Pos_232;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_232 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_232;   
  
  Energy_Bin_Pos_233 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_233   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_233 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E233_C1_L_Pos and PEAK_C1_Pos <= s_E233_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_233 <= s_Energy_Bin_Pos_233 +'1';
		 Energy_Bin_Pos_Rdy_233 <= '1';
		else
		 s_Energy_Bin_Pos_233 <= s_Energy_Bin_Pos_233;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_233 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_233;   
  
  Energy_Bin_Pos_234 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_234   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_234 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E234_C1_L_Pos and PEAK_C1_Pos <= s_E234_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_234 <= s_Energy_Bin_Pos_234 +'1';
		 Energy_Bin_Pos_Rdy_234 <= '1';
		else
		 s_Energy_Bin_Pos_234 <= s_Energy_Bin_Pos_234;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_234 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_234;   
 
 
  Energy_Bin_Pos_235 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_235   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_235 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E235_C1_L_Pos and PEAK_C1_Pos <= s_E235_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_235 <= s_Energy_Bin_Pos_235 +'1';
		 Energy_Bin_Pos_Rdy_235 <= '1';
		else
		 s_Energy_Bin_Pos_235 <= s_Energy_Bin_Pos_235;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_235 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_235;  
 
  
  Energy_Bin_Pos_236 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_236   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_236 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E236_C1_L_Pos and PEAK_C1_Pos <= s_E236_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_236 <= s_Energy_Bin_Pos_236 +'1';
		 Energy_Bin_Pos_Rdy_236 <= '1';
		else
		 s_Energy_Bin_Pos_236 <= s_Energy_Bin_Pos_236;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_236 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_236;   
  
 Energy_Bin_Pos_237 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_237   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_237 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E237_C1_L_Pos and PEAK_C1_Pos <= s_E237_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_237 <= s_Energy_Bin_Pos_237 +'1';
		 Energy_Bin_Pos_Rdy_237 <= '1';
		else
		 s_Energy_Bin_Pos_237 <= s_Energy_Bin_Pos_237;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_237 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_237;   
  
  Energy_Bin_Pos_238 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_238   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_238 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E238_C1_L_Pos and PEAK_C1_Pos <= s_E238_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_238 <= s_Energy_Bin_Pos_238 +'1';
		 Energy_Bin_Pos_Rdy_238 <= '1';
		else
		 s_Energy_Bin_Pos_238 <= s_Energy_Bin_Pos_238;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_238 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_238;   
  
  Energy_Bin_Pos_239 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_239   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_239 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E239_C1_L_Pos and PEAK_C1_Pos <= s_E239_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_239 <= s_Energy_Bin_Pos_239 +'1';
		 Energy_Bin_Pos_Rdy_239 <= '1';
		else
		 s_Energy_Bin_Pos_239 <= s_Energy_Bin_Pos_239;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_239 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_239;         
  
     Energy_Bin_Pos_240 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_240   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_240 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E240_C1_L_Pos and PEAK_C1_Pos <= s_E240_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_240 <= s_Energy_Bin_Pos_240 +'1';
		 Energy_Bin_Pos_Rdy_240 <= '1';
		else
		 s_Energy_Bin_Pos_240 <= s_Energy_Bin_Pos_240;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_240 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_240;    
  
  Energy_Bin_Pos_241 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_241   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_241 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E241_C1_L_Pos and PEAK_C1_Pos <= s_E241_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_241 <= s_Energy_Bin_Pos_241 +'1';
		 Energy_Bin_Pos_Rdy_241 <= '1';
		else
		 s_Energy_Bin_Pos_241 <= s_Energy_Bin_Pos_241;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_241 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_241;   
  
  Energy_Bin_Pos_242 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_242   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_242 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E242_C1_L_Pos and PEAK_C1_Pos <= s_E242_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_242 <= s_Energy_Bin_Pos_242 +'1';
		 Energy_Bin_Pos_Rdy_242 <= '1';
		else
		 s_Energy_Bin_Pos_242 <= s_Energy_Bin_Pos_242;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_242 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_242;   
  
  Energy_Bin_Pos_243 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_243   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_243 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E243_C1_L_Pos and PEAK_C1_Pos <= s_E243_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_243 <= s_Energy_Bin_Pos_243 +'1';
		 Energy_Bin_Pos_Rdy_243 <= '1';
		else
		 s_Energy_Bin_Pos_243 <= s_Energy_Bin_Pos_243;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_243 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_243;   
  
  Energy_Bin_Pos_244 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_244   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_244 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E244_C1_L_Pos and PEAK_C1_Pos <= s_E244_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_244 <= s_Energy_Bin_Pos_244 +'1';
		 Energy_Bin_Pos_Rdy_244 <= '1';
		else
		 s_Energy_Bin_Pos_244 <= s_Energy_Bin_Pos_244;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_244 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_244;   
 
 
  Energy_Bin_Pos_245 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_245   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_245 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E245_C1_L_Pos and PEAK_C1_Pos <= s_E245_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_245 <= s_Energy_Bin_Pos_245 +'1';
		 Energy_Bin_Pos_Rdy_245 <= '1';
		else
		 s_Energy_Bin_Pos_245 <= s_Energy_Bin_Pos_245;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_245 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_245;  
 
  
  Energy_Bin_Pos_246 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_246   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_246 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E246_C1_L_Pos and PEAK_C1_Pos <= s_E246_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_246 <= s_Energy_Bin_Pos_246 +'1';
		 Energy_Bin_Pos_Rdy_246 <= '1';
		else
		 s_Energy_Bin_Pos_246 <= s_Energy_Bin_Pos_246;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_246 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_246;   
  
 Energy_Bin_Pos_247 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_247   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_247 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E247_C1_L_Pos and PEAK_C1_Pos <= s_E247_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_247 <= s_Energy_Bin_Pos_247 +'1';
		 Energy_Bin_Pos_Rdy_247 <= '1';
		else
		 s_Energy_Bin_Pos_247 <= s_Energy_Bin_Pos_247;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_247 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_247;   
  
  Energy_Bin_Pos_248 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_248   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_248 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E248_C1_L_Pos and PEAK_C1_Pos <= s_E248_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_248 <= s_Energy_Bin_Pos_248 +'1';
		 Energy_Bin_Pos_Rdy_248 <= '1';
		else
		 s_Energy_Bin_Pos_248 <= s_Energy_Bin_Pos_248;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_248 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_248;   
  
  Energy_Bin_Pos_249 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_249   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_249 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E249_C1_L_Pos and PEAK_C1_Pos <= s_E249_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_249 <= s_Energy_Bin_Pos_249 +'1';
		 Energy_Bin_Pos_Rdy_249 <= '1';
		else
		 s_Energy_Bin_Pos_249 <= s_Energy_Bin_Pos_249;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_249 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_249;          
  
  
     Energy_Bin_Pos_250 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_250   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_250 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E250_C1_L_Pos and PEAK_C1_Pos <= s_E250_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_250 <= s_Energy_Bin_Pos_250 +'1';
		 Energy_Bin_Pos_Rdy_250 <= '1';
		else
		 s_Energy_Bin_Pos_250 <= s_Energy_Bin_Pos_250;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_250 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_250;    
  
  Energy_Bin_Pos_251 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_251   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_251 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E251_C1_L_Pos and PEAK_C1_Pos <= s_E251_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_251 <= s_Energy_Bin_Pos_251 +'1';
		 Energy_Bin_Pos_Rdy_251 <= '1';
		else
		 s_Energy_Bin_Pos_251 <= s_Energy_Bin_Pos_251;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_251 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_251;   
  
  Energy_Bin_Pos_252 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_252   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_252 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E252_C1_L_Pos and PEAK_C1_Pos <= s_E252_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_252 <= s_Energy_Bin_Pos_252 +'1';
		 Energy_Bin_Pos_Rdy_252 <= '1';
		else
		 s_Energy_Bin_Pos_252 <= s_Energy_Bin_Pos_252;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_252 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_252;   
  
  Energy_Bin_Pos_253 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_253   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_253 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E253_C1_L_Pos and PEAK_C1_Pos <= s_E253_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_253 <= s_Energy_Bin_Pos_253 +'1';
		 Energy_Bin_Pos_Rdy_253 <= '1';
		else
		 s_Energy_Bin_Pos_253 <= s_Energy_Bin_Pos_253;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_253 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_253;   
  
  Energy_Bin_Pos_254 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_254   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_254 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E254_C1_L_Pos and PEAK_C1_Pos <= s_E254_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_254 <= s_Energy_Bin_Pos_254 +'1';
		 Energy_Bin_Pos_Rdy_254 <= '1';
		else
		 s_Energy_Bin_Pos_254 <= s_Energy_Bin_Pos_254;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_254 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_254;   
 
 
  Energy_Bin_Pos_255 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_255   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_255 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E255_C1_L_Pos and PEAK_C1_Pos <= s_E255_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_255 <= s_Energy_Bin_Pos_255 +'1';
		 Energy_Bin_Pos_Rdy_255 <= '1';
		else
		 s_Energy_Bin_Pos_255 <= s_Energy_Bin_Pos_255;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_255 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_255;  
 
  
  Energy_Bin_Pos_256 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_256   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_256 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E256_C1_L_Pos and PEAK_C1_Pos <= s_E256_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_256 <= s_Energy_Bin_Pos_256 +'1';
		 Energy_Bin_Pos_Rdy_256 <= '1';
		else
		 s_Energy_Bin_Pos_256 <= s_Energy_Bin_Pos_256;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_256 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_256;   
  
 Energy_Bin_Pos_257 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_257   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_257 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E257_C1_L_Pos and PEAK_C1_Pos <= s_E257_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_257 <= s_Energy_Bin_Pos_257 +'1';
		 Energy_Bin_Pos_Rdy_257 <= '1';
		else
		 s_Energy_Bin_Pos_257 <= s_Energy_Bin_Pos_257;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_257 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_257;   
  
  Energy_Bin_Pos_258 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_258   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_258 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E258_C1_L_Pos and PEAK_C1_Pos <= s_E258_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_258 <= s_Energy_Bin_Pos_258 +'1';
		 Energy_Bin_Pos_Rdy_258 <= '1';
		else
		 s_Energy_Bin_Pos_258 <= s_Energy_Bin_Pos_258;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_258 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_258;   
  
  Energy_Bin_Pos_259 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_259   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_259 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E259_C1_L_Pos and PEAK_C1_Pos <= s_E259_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_259 <= s_Energy_Bin_Pos_259 +'1';
		 Energy_Bin_Pos_Rdy_259 <= '1';
		else
		 s_Energy_Bin_Pos_259 <= s_Energy_Bin_Pos_259;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_259 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_259;           
  
     Energy_Bin_Pos_260 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_260   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_260 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E260_C1_L_Pos and PEAK_C1_Pos <= s_E260_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_260 <= s_Energy_Bin_Pos_260 +'1';
		 Energy_Bin_Pos_Rdy_260 <= '1';
		else
		 s_Energy_Bin_Pos_260 <= s_Energy_Bin_Pos_260;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_260 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_260;    
  
  Energy_Bin_Pos_261 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_261   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_261 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E261_C1_L_Pos and PEAK_C1_Pos <= s_E261_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_261 <= s_Energy_Bin_Pos_261 +'1';
		 Energy_Bin_Pos_Rdy_261 <= '1';
		else
		 s_Energy_Bin_Pos_261 <= s_Energy_Bin_Pos_261;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_261 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_261;   
  
  Energy_Bin_Pos_262 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_262   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_262 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E262_C1_L_Pos and PEAK_C1_Pos <= s_E262_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_262 <= s_Energy_Bin_Pos_262 +'1';
		 Energy_Bin_Pos_Rdy_262 <= '1';
		else
		 s_Energy_Bin_Pos_262 <= s_Energy_Bin_Pos_262;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_262 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_262;   
  
  Energy_Bin_Pos_263 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_263   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_263 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E263_C1_L_Pos and PEAK_C1_Pos <= s_E263_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_263 <= s_Energy_Bin_Pos_263 +'1';
		 Energy_Bin_Pos_Rdy_263 <= '1';
		else
		 s_Energy_Bin_Pos_263 <= s_Energy_Bin_Pos_263;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_263 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_263;   
  
  Energy_Bin_Pos_264 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_264   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_264 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E264_C1_L_Pos and PEAK_C1_Pos <= s_E264_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_264 <= s_Energy_Bin_Pos_264 +'1';
		 Energy_Bin_Pos_Rdy_264 <= '1';
		else
		 s_Energy_Bin_Pos_264 <= s_Energy_Bin_Pos_264;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_264 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_264;   
 
 
  Energy_Bin_Pos_265 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_265   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_265 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E265_C1_L_Pos and PEAK_C1_Pos <= s_E265_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_265 <= s_Energy_Bin_Pos_265 +'1';
		 Energy_Bin_Pos_Rdy_265 <= '1';
		else
		 s_Energy_Bin_Pos_265 <= s_Energy_Bin_Pos_265;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_265 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_265;  
 
  
  Energy_Bin_Pos_266 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_266   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_266 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E266_C1_L_Pos and PEAK_C1_Pos <= s_E266_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_266 <= s_Energy_Bin_Pos_266 +'1';
		 Energy_Bin_Pos_Rdy_266 <= '1';
		else
		 s_Energy_Bin_Pos_266 <= s_Energy_Bin_Pos_266;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_266 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_266;   
  
 Energy_Bin_Pos_267 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_267   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_267 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E267_C1_L_Pos and PEAK_C1_Pos <= s_E267_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_267 <= s_Energy_Bin_Pos_267 +'1';
		 Energy_Bin_Pos_Rdy_267 <= '1';
		else
		 s_Energy_Bin_Pos_267 <= s_Energy_Bin_Pos_267;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_267 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_267;   
  
  Energy_Bin_Pos_268 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_268   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_268 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E268_C1_L_Pos and PEAK_C1_Pos <= s_E268_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_268 <= s_Energy_Bin_Pos_268 +'1';
		 Energy_Bin_Pos_Rdy_268 <= '1';
		else
		 s_Energy_Bin_Pos_268 <= s_Energy_Bin_Pos_268;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_268 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_268;   
  
  Energy_Bin_Pos_269 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_269   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_269 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E269_C1_L_Pos and PEAK_C1_Pos <= s_E269_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_269 <= s_Energy_Bin_Pos_269 +'1';
		 Energy_Bin_Pos_Rdy_269 <= '1';
		else
		 s_Energy_Bin_Pos_269 <= s_Energy_Bin_Pos_269;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_269 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_269;         
  
     Energy_Bin_Pos_270 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_270   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_270 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E270_C1_L_Pos and PEAK_C1_Pos <= s_E270_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_270 <= s_Energy_Bin_Pos_270 +'1';
		 Energy_Bin_Pos_Rdy_270 <= '1';
		else
		 s_Energy_Bin_Pos_270 <= s_Energy_Bin_Pos_270;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_270 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_270;    
  
  Energy_Bin_Pos_271 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_271   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_271 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E271_C1_L_Pos and PEAK_C1_Pos <= s_E271_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_271 <= s_Energy_Bin_Pos_271 +'1';
		 Energy_Bin_Pos_Rdy_271 <= '1';
		else
		 s_Energy_Bin_Pos_271 <= s_Energy_Bin_Pos_271;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_271 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_271;   
  
  Energy_Bin_Pos_272 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_272   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_272 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E272_C1_L_Pos and PEAK_C1_Pos <= s_E272_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_272 <= s_Energy_Bin_Pos_272 +'1';
		 Energy_Bin_Pos_Rdy_272 <= '1';
		else
		 s_Energy_Bin_Pos_272 <= s_Energy_Bin_Pos_272;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_272 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_272;   
  
  Energy_Bin_Pos_273 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_273   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_273 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E273_C1_L_Pos and PEAK_C1_Pos <= s_E273_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_273 <= s_Energy_Bin_Pos_273 +'1';
		 Energy_Bin_Pos_Rdy_273 <= '1';
		else
		 s_Energy_Bin_Pos_273 <= s_Energy_Bin_Pos_273;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_273 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_273;   
  
  Energy_Bin_Pos_274 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_274   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_274 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E274_C1_L_Pos and PEAK_C1_Pos <= s_E274_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_274 <= s_Energy_Bin_Pos_274 +'1';
		 Energy_Bin_Pos_Rdy_274 <= '1';
		else
		 s_Energy_Bin_Pos_274 <= s_Energy_Bin_Pos_274;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_274 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_274;   
 
 
  Energy_Bin_Pos_275 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_275   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_275 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E275_C1_L_Pos and PEAK_C1_Pos <= s_E275_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_275 <= s_Energy_Bin_Pos_275 +'1';
		 Energy_Bin_Pos_Rdy_275 <= '1';
		else
		 s_Energy_Bin_Pos_275 <= s_Energy_Bin_Pos_275;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_275 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_275;  
 
  
  Energy_Bin_Pos_276 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_276   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_276 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E276_C1_L_Pos and PEAK_C1_Pos <= s_E276_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_276 <= s_Energy_Bin_Pos_276 +'1';
		 Energy_Bin_Pos_Rdy_276 <= '1';
		else
		 s_Energy_Bin_Pos_276 <= s_Energy_Bin_Pos_276;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_276 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_276;   
  
 Energy_Bin_Pos_277 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_277   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_277 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E277_C1_L_Pos and PEAK_C1_Pos <= s_E277_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_277 <= s_Energy_Bin_Pos_277 +'1';
		 Energy_Bin_Pos_Rdy_277 <= '1';
		else
		 s_Energy_Bin_Pos_277 <= s_Energy_Bin_Pos_277;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_277 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_277;   
  
  Energy_Bin_Pos_278 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_278   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_278 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E278_C1_L_Pos and PEAK_C1_Pos <= s_E278_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_278 <= s_Energy_Bin_Pos_278 +'1';
		 Energy_Bin_Pos_Rdy_278 <= '1';
		else
		 s_Energy_Bin_Pos_278 <= s_Energy_Bin_Pos_278;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_278 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_278;   
  
  Energy_Bin_Pos_279 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_279   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_279 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E279_C1_L_Pos and PEAK_C1_Pos <= s_E279_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_279 <= s_Energy_Bin_Pos_279 +'1';
		 Energy_Bin_Pos_Rdy_279 <= '1';
		else
		 s_Energy_Bin_Pos_279 <= s_Energy_Bin_Pos_279;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_279 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_279;       
  
     Energy_Bin_Pos_280 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_280   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_280 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E280_C1_L_Pos and PEAK_C1_Pos <= s_E280_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_280 <= s_Energy_Bin_Pos_280 +'1';
		 Energy_Bin_Pos_Rdy_280 <= '1';
		else
		 s_Energy_Bin_Pos_280 <= s_Energy_Bin_Pos_280;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_280 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_280;    
  
  Energy_Bin_Pos_281 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_281   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_281 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E281_C1_L_Pos and PEAK_C1_Pos <= s_E281_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_281 <= s_Energy_Bin_Pos_281 +'1';
		 Energy_Bin_Pos_Rdy_281 <= '1';
		else
		 s_Energy_Bin_Pos_281 <= s_Energy_Bin_Pos_281;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_281 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_281;   
  
  Energy_Bin_Pos_282 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_282   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_282 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E282_C1_L_Pos and PEAK_C1_Pos <= s_E282_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_282 <= s_Energy_Bin_Pos_282 +'1';
		 Energy_Bin_Pos_Rdy_282 <= '1';
		else
		 s_Energy_Bin_Pos_282 <= s_Energy_Bin_Pos_282;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_282 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_282;   
  
  Energy_Bin_Pos_283 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_283   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_283 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E283_C1_L_Pos and PEAK_C1_Pos <= s_E283_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_283 <= s_Energy_Bin_Pos_283 +'1';
		 Energy_Bin_Pos_Rdy_283 <= '1';
		else
		 s_Energy_Bin_Pos_283 <= s_Energy_Bin_Pos_283;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_283 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_283;   
  
  Energy_Bin_Pos_284 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_284   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_284 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E284_C1_L_Pos and PEAK_C1_Pos <= s_E284_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_284 <= s_Energy_Bin_Pos_284 +'1';
		 Energy_Bin_Pos_Rdy_284 <= '1';
		else
		 s_Energy_Bin_Pos_284 <= s_Energy_Bin_Pos_284;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_284 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_284;   
 
 
  Energy_Bin_Pos_285 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_285   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_285 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E285_C1_L_Pos and PEAK_C1_Pos <= s_E285_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_285 <= s_Energy_Bin_Pos_285 +'1';
		 Energy_Bin_Pos_Rdy_285 <= '1';
		else
		 s_Energy_Bin_Pos_285 <= s_Energy_Bin_Pos_285;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_285 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_285;  
 
  
  Energy_Bin_Pos_286 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_286   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_286 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E286_C1_L_Pos and PEAK_C1_Pos <= s_E286_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_286 <= s_Energy_Bin_Pos_286 +'1';
		 Energy_Bin_Pos_Rdy_286 <= '1';
		else
		 s_Energy_Bin_Pos_286 <= s_Energy_Bin_Pos_286;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_286 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_286;   
  
 Energy_Bin_Pos_287 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_287   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_287 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E287_C1_L_Pos and PEAK_C1_Pos <= s_E287_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_287 <= s_Energy_Bin_Pos_287 +'1';
		 Energy_Bin_Pos_Rdy_287 <= '1';
		else
		 s_Energy_Bin_Pos_287 <= s_Energy_Bin_Pos_287;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_287 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_287;   
  
  Energy_Bin_Pos_288 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_288   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_288 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E288_C1_L_Pos and PEAK_C1_Pos <= s_E288_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_288 <= s_Energy_Bin_Pos_288 +'1';
		 Energy_Bin_Pos_Rdy_288 <= '1';
		else
		 s_Energy_Bin_Pos_288 <= s_Energy_Bin_Pos_288;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_288 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_288;   
  
  Energy_Bin_Pos_289 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_289   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_289 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E289_C1_L_Pos and PEAK_C1_Pos <= s_E289_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_289 <= s_Energy_Bin_Pos_289 +'1';
		 Energy_Bin_Pos_Rdy_289 <= '1';
		else
		 s_Energy_Bin_Pos_289 <= s_Energy_Bin_Pos_289;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_289 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_289;      
  
     Energy_Bin_Pos_290 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_290   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_290 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E290_C1_L_Pos and PEAK_C1_Pos <= s_E290_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_290 <= s_Energy_Bin_Pos_290 +'1';
		 Energy_Bin_Pos_Rdy_290 <= '1';
		else
		 s_Energy_Bin_Pos_290 <= s_Energy_Bin_Pos_290;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_290 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_290;    
  
  Energy_Bin_Pos_291 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_291   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_291 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E291_C1_L_Pos and PEAK_C1_Pos <= s_E291_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_291 <= s_Energy_Bin_Pos_291 +'1';
		 Energy_Bin_Pos_Rdy_291 <= '1';
		else
		 s_Energy_Bin_Pos_291 <= s_Energy_Bin_Pos_291;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_291 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_291;   
  
  Energy_Bin_Pos_292 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_292   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_292 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E292_C1_L_Pos and PEAK_C1_Pos <= s_E292_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_292 <= s_Energy_Bin_Pos_292 +'1';
		 Energy_Bin_Pos_Rdy_292 <= '1';
		else
		 s_Energy_Bin_Pos_292 <= s_Energy_Bin_Pos_292;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_292 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_292;   
  
  Energy_Bin_Pos_293 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_293   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_293 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E293_C1_L_Pos and PEAK_C1_Pos <= s_E293_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_293 <= s_Energy_Bin_Pos_293 +'1';
		 Energy_Bin_Pos_Rdy_293 <= '1';
		else
		 s_Energy_Bin_Pos_293 <= s_Energy_Bin_Pos_293;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_293 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_293;   
  
  Energy_Bin_Pos_294 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_294   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_294 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E294_C1_L_Pos and PEAK_C1_Pos <= s_E294_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_294 <= s_Energy_Bin_Pos_294 +'1';
		 Energy_Bin_Pos_Rdy_294 <= '1';
		else
		 s_Energy_Bin_Pos_294 <= s_Energy_Bin_Pos_294;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_294 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_294;   
 
 
  Energy_Bin_Pos_295 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_295   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_295 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E295_C1_L_Pos and PEAK_C1_Pos <= s_E295_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_295 <= s_Energy_Bin_Pos_295 +'1';
		 Energy_Bin_Pos_Rdy_295 <= '1';
		else
		 s_Energy_Bin_Pos_295 <= s_Energy_Bin_Pos_295;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_295 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_295;  
 
  
  Energy_Bin_Pos_296 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_296   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_296 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E296_C1_L_Pos and PEAK_C1_Pos <= s_E296_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_296 <= s_Energy_Bin_Pos_296 +'1';
		 Energy_Bin_Pos_Rdy_296 <= '1';
		else
		 s_Energy_Bin_Pos_296 <= s_Energy_Bin_Pos_296;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_296 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_296;   
  
 Energy_Bin_Pos_297 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_297   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_297 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E297_C1_L_Pos and PEAK_C1_Pos <= s_E297_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_297 <= s_Energy_Bin_Pos_297 +'1';
		 Energy_Bin_Pos_Rdy_297 <= '1';
		else
		 s_Energy_Bin_Pos_297 <= s_Energy_Bin_Pos_297;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_297 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_297;   
  
  Energy_Bin_Pos_298 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_298   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_298 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E298_C1_L_Pos and PEAK_C1_Pos <= s_E298_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_298 <= s_Energy_Bin_Pos_298 +'1';
		 Energy_Bin_Pos_Rdy_298 <= '1';
		else
		 s_Energy_Bin_Pos_298 <= s_Energy_Bin_Pos_298;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_298 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_298;   
  
  Energy_Bin_Pos_299 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_299   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_299 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E299_C1_L_Pos and PEAK_C1_Pos <= s_E299_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_299 <= s_Energy_Bin_Pos_299 +'1';
		 Energy_Bin_Pos_Rdy_299 <= '1';
		else
		 s_Energy_Bin_Pos_299 <= s_Energy_Bin_Pos_299;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_299 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_299;      

     Energy_Bin_Pos_300 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_300   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_300 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E300_C1_L_Pos and PEAK_C1_Pos <= s_E300_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_300 <= s_Energy_Bin_Pos_300 +'1';
		 Energy_Bin_Pos_Rdy_300 <= '1';
		else
		 s_Energy_Bin_Pos_300 <= s_Energy_Bin_Pos_300;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_300 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_300;    
  
  Energy_Bin_Pos_301 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_301   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_301 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E301_C1_L_Pos and PEAK_C1_Pos <= s_E301_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_301 <= s_Energy_Bin_Pos_301 +'1';
		 Energy_Bin_Pos_Rdy_301 <= '1';
		else
		 s_Energy_Bin_Pos_301 <= s_Energy_Bin_Pos_301;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_301 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_301;   
  
  Energy_Bin_Pos_302 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_302   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_302 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E302_C1_L_Pos and PEAK_C1_Pos <= s_E302_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_302 <= s_Energy_Bin_Pos_302 +'1';
		 Energy_Bin_Pos_Rdy_302 <= '1';
		else
		 s_Energy_Bin_Pos_302 <= s_Energy_Bin_Pos_302;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_302 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_302;   
  
  Energy_Bin_Pos_303 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_303   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_303 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E303_C1_L_Pos and PEAK_C1_Pos <= s_E303_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_303 <= s_Energy_Bin_Pos_303 +'1';
		 Energy_Bin_Pos_Rdy_303 <= '1';
		else
		 s_Energy_Bin_Pos_303 <= s_Energy_Bin_Pos_303;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_303 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_303;   
  
  Energy_Bin_Pos_304 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_304   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_304 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E304_C1_L_Pos and PEAK_C1_Pos <= s_E304_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_304 <= s_Energy_Bin_Pos_304 +'1';
		 Energy_Bin_Pos_Rdy_304 <= '1';
		else
		 s_Energy_Bin_Pos_304 <= s_Energy_Bin_Pos_304;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_304 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_304;   
 
 
  Energy_Bin_Pos_305 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_305   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_305 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E305_C1_L_Pos and PEAK_C1_Pos <= s_E305_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_305 <= s_Energy_Bin_Pos_305 +'1';
		 Energy_Bin_Pos_Rdy_305 <= '1';
		else
		 s_Energy_Bin_Pos_305 <= s_Energy_Bin_Pos_305;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_305 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_305;  
 
  
  Energy_Bin_Pos_306 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_306   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_306 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E306_C1_L_Pos and PEAK_C1_Pos <= s_E306_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_306 <= s_Energy_Bin_Pos_306 +'1';
		 Energy_Bin_Pos_Rdy_306 <= '1';
		else
		 s_Energy_Bin_Pos_306 <= s_Energy_Bin_Pos_306;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_306 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_306;   
  
 Energy_Bin_Pos_307 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_307   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_307 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E307_C1_L_Pos and PEAK_C1_Pos <= s_E307_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_307 <= s_Energy_Bin_Pos_307 +'1';
		 Energy_Bin_Pos_Rdy_307 <= '1';
		else
		 s_Energy_Bin_Pos_307 <= s_Energy_Bin_Pos_307;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_307 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_307;   
  
  Energy_Bin_Pos_308 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_308   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_308 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E308_C1_L_Pos and PEAK_C1_Pos <= s_E308_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_308 <= s_Energy_Bin_Pos_308 +'1';
		 Energy_Bin_Pos_Rdy_308 <= '1';
		else
		 s_Energy_Bin_Pos_308 <= s_Energy_Bin_Pos_308;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_308 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_308;   
  
  Energy_Bin_Pos_309 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_309   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_309 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E309_C1_L_Pos and PEAK_C1_Pos <= s_E309_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_309 <= s_Energy_Bin_Pos_309 +'1';
		 Energy_Bin_Pos_Rdy_309 <= '1';
		else
		 s_Energy_Bin_Pos_309 <= s_Energy_Bin_Pos_309;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_309 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_309;      
  
     Energy_Bin_Pos_310 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_310   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_310 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E310_C1_L_Pos and PEAK_C1_Pos <= s_E310_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_310 <= s_Energy_Bin_Pos_310 +'1';
		 Energy_Bin_Pos_Rdy_310 <= '1';
		else
		 s_Energy_Bin_Pos_310 <= s_Energy_Bin_Pos_310;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_310 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_310;    
  
  Energy_Bin_Pos_311 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_311   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_311 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E311_C1_L_Pos and PEAK_C1_Pos <= s_E311_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_311 <= s_Energy_Bin_Pos_311 +'1';
		 Energy_Bin_Pos_Rdy_311 <= '1';
		else
		 s_Energy_Bin_Pos_311 <= s_Energy_Bin_Pos_311;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_311 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_311;   
  
  Energy_Bin_Pos_312 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_312   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_312 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E312_C1_L_Pos and PEAK_C1_Pos <= s_E312_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_312 <= s_Energy_Bin_Pos_312 +'1';
		 Energy_Bin_Pos_Rdy_312 <= '1';
		else
		 s_Energy_Bin_Pos_312 <= s_Energy_Bin_Pos_312;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_312 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_312;   
  
  Energy_Bin_Pos_313 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_313   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_313 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E313_C1_L_Pos and PEAK_C1_Pos <= s_E313_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_313 <= s_Energy_Bin_Pos_313 +'1';
		 Energy_Bin_Pos_Rdy_313 <= '1';
		else
		 s_Energy_Bin_Pos_313 <= s_Energy_Bin_Pos_313;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_313 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_313;   
  
  Energy_Bin_Pos_314 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_314   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_314 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E314_C1_L_Pos and PEAK_C1_Pos <= s_E314_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_314 <= s_Energy_Bin_Pos_314 +'1';
		 Energy_Bin_Pos_Rdy_314 <= '1';
		else
		 s_Energy_Bin_Pos_314 <= s_Energy_Bin_Pos_314;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_314 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_314;   
 
 
  Energy_Bin_Pos_315 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_315   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_315 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E315_C1_L_Pos and PEAK_C1_Pos <= s_E315_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_315 <= s_Energy_Bin_Pos_315 +'1';
		 Energy_Bin_Pos_Rdy_315 <= '1';
		else
		 s_Energy_Bin_Pos_315 <= s_Energy_Bin_Pos_315;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_315 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_315;  
 
  
  Energy_Bin_Pos_316 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_316   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_316 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E316_C1_L_Pos and PEAK_C1_Pos <= s_E316_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_316 <= s_Energy_Bin_Pos_316 +'1';
		 Energy_Bin_Pos_Rdy_316 <= '1';
		else
		 s_Energy_Bin_Pos_316 <= s_Energy_Bin_Pos_316;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_316 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_316;   
  
 Energy_Bin_Pos_317 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_317   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_317 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E317_C1_L_Pos and PEAK_C1_Pos <= s_E317_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_317 <= s_Energy_Bin_Pos_317 +'1';
		 Energy_Bin_Pos_Rdy_317 <= '1';
		else
		 s_Energy_Bin_Pos_317 <= s_Energy_Bin_Pos_317;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_317 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_317;   
  
  Energy_Bin_Pos_318 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_318   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_318 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E318_C1_L_Pos and PEAK_C1_Pos <= s_E318_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_318 <= s_Energy_Bin_Pos_318 +'1';
		 Energy_Bin_Pos_Rdy_318 <= '1';
		else
		 s_Energy_Bin_Pos_318 <= s_Energy_Bin_Pos_318;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_318 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_318;   
  
  Energy_Bin_Pos_319 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_319   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_319 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E319_C1_L_Pos and PEAK_C1_Pos <= s_E319_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_319 <= s_Energy_Bin_Pos_319 +'1';
		 Energy_Bin_Pos_Rdy_319 <= '1';
		else
		 s_Energy_Bin_Pos_319 <= s_Energy_Bin_Pos_319;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_319 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_319;       
  
     Energy_Bin_Pos_320 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_320   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_320 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E320_C1_L_Pos and PEAK_C1_Pos <= s_E320_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_320 <= s_Energy_Bin_Pos_320 +'1';
		 Energy_Bin_Pos_Rdy_320 <= '1';
		else
		 s_Energy_Bin_Pos_320 <= s_Energy_Bin_Pos_320;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_320 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_320;    
  
  Energy_Bin_Pos_321 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_321   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_321 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E321_C1_L_Pos and PEAK_C1_Pos <= s_E321_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_321 <= s_Energy_Bin_Pos_321 +'1';
		 Energy_Bin_Pos_Rdy_321 <= '1';
		else
		 s_Energy_Bin_Pos_321 <= s_Energy_Bin_Pos_321;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_321 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_321;   
  
  Energy_Bin_Pos_322 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_322   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_322 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E322_C1_L_Pos and PEAK_C1_Pos <= s_E322_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_322 <= s_Energy_Bin_Pos_322 +'1';
		 Energy_Bin_Pos_Rdy_322 <= '1';
		else
		 s_Energy_Bin_Pos_322 <= s_Energy_Bin_Pos_322;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_322 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_322;   
  
  Energy_Bin_Pos_323 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_323   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_323 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E323_C1_L_Pos and PEAK_C1_Pos <= s_E323_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_323 <= s_Energy_Bin_Pos_323 +'1';
		 Energy_Bin_Pos_Rdy_323 <= '1';
		else
		 s_Energy_Bin_Pos_323 <= s_Energy_Bin_Pos_323;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_323 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_323;   
  
  Energy_Bin_Pos_324 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_324   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_324 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E324_C1_L_Pos and PEAK_C1_Pos <= s_E324_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_324 <= s_Energy_Bin_Pos_324 +'1';
		 Energy_Bin_Pos_Rdy_324 <= '1';
		else
		 s_Energy_Bin_Pos_324 <= s_Energy_Bin_Pos_324;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_324 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_324;   
 
 
  Energy_Bin_Pos_325 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_325   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_325 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E325_C1_L_Pos and PEAK_C1_Pos <= s_E325_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_325 <= s_Energy_Bin_Pos_325 +'1';
		 Energy_Bin_Pos_Rdy_325 <= '1';
		else
		 s_Energy_Bin_Pos_325 <= s_Energy_Bin_Pos_325;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_325 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_325;  
 
  
  Energy_Bin_Pos_326 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_326   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_326 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E326_C1_L_Pos and PEAK_C1_Pos <= s_E326_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_326 <= s_Energy_Bin_Pos_326 +'1';
		 Energy_Bin_Pos_Rdy_326 <= '1';
		else
		 s_Energy_Bin_Pos_326 <= s_Energy_Bin_Pos_326;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_326 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_326;   
  
 Energy_Bin_Pos_327 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_327   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_327 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E327_C1_L_Pos and PEAK_C1_Pos <= s_E327_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_327 <= s_Energy_Bin_Pos_327 +'1';
		 Energy_Bin_Pos_Rdy_327 <= '1';
		else
		 s_Energy_Bin_Pos_327 <= s_Energy_Bin_Pos_327;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_327 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_327;   
  
  Energy_Bin_Pos_328 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_328   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_328 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E328_C1_L_Pos and PEAK_C1_Pos <= s_E328_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_328 <= s_Energy_Bin_Pos_328 +'1';
		 Energy_Bin_Pos_Rdy_328 <= '1';
		else
		 s_Energy_Bin_Pos_328 <= s_Energy_Bin_Pos_328;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_328 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_328;   
  
  Energy_Bin_Pos_329 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_329   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_329 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E329_C1_L_Pos and PEAK_C1_Pos <= s_E329_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_329 <= s_Energy_Bin_Pos_329 +'1';
		 Energy_Bin_Pos_Rdy_329 <= '1';
		else
		 s_Energy_Bin_Pos_329 <= s_Energy_Bin_Pos_329;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_329 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_329;        
  
     Energy_Bin_Pos_330 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_330   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_330 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E330_C1_L_Pos and PEAK_C1_Pos <= s_E330_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_330 <= s_Energy_Bin_Pos_330 +'1';
		 Energy_Bin_Pos_Rdy_330 <= '1';
		else
		 s_Energy_Bin_Pos_330 <= s_Energy_Bin_Pos_330;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_330 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_330;    
  
  Energy_Bin_Pos_331 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_331   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_331 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E331_C1_L_Pos and PEAK_C1_Pos <= s_E331_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_331 <= s_Energy_Bin_Pos_331 +'1';
		 Energy_Bin_Pos_Rdy_331 <= '1';
		else
		 s_Energy_Bin_Pos_331 <= s_Energy_Bin_Pos_331;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_331 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_331;   
  
  Energy_Bin_Pos_332 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_332   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_332 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E332_C1_L_Pos and PEAK_C1_Pos <= s_E332_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_332 <= s_Energy_Bin_Pos_332 +'1';
		 Energy_Bin_Pos_Rdy_332 <= '1';
		else
		 s_Energy_Bin_Pos_332 <= s_Energy_Bin_Pos_332;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_332 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_332;   
  
  Energy_Bin_Pos_333 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_333   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_333 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E333_C1_L_Pos and PEAK_C1_Pos <= s_E333_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_333 <= s_Energy_Bin_Pos_333 +'1';
		 Energy_Bin_Pos_Rdy_333 <= '1';
		else
		 s_Energy_Bin_Pos_333 <= s_Energy_Bin_Pos_333;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_333 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_333;   
  
  Energy_Bin_Pos_334 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_334   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_334 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E334_C1_L_Pos and PEAK_C1_Pos <= s_E334_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_334 <= s_Energy_Bin_Pos_334 +'1';
		 Energy_Bin_Pos_Rdy_334 <= '1';
		else
		 s_Energy_Bin_Pos_334 <= s_Energy_Bin_Pos_334;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_334 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_334;   
 
 
  Energy_Bin_Pos_335 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_335   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_335 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E335_C1_L_Pos and PEAK_C1_Pos <= s_E335_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_335 <= s_Energy_Bin_Pos_335 +'1';
		 Energy_Bin_Pos_Rdy_335 <= '1';
		else
		 s_Energy_Bin_Pos_335 <= s_Energy_Bin_Pos_335;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_335 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_335;  
 
  
  Energy_Bin_Pos_336 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_336   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_336 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E336_C1_L_Pos and PEAK_C1_Pos <= s_E336_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_336 <= s_Energy_Bin_Pos_336 +'1';
		 Energy_Bin_Pos_Rdy_336 <= '1';
		else
		 s_Energy_Bin_Pos_336 <= s_Energy_Bin_Pos_336;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_336 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_336;   
  
 Energy_Bin_Pos_337 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_337   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_337 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E337_C1_L_Pos and PEAK_C1_Pos <= s_E337_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_337 <= s_Energy_Bin_Pos_337 +'1';
		 Energy_Bin_Pos_Rdy_337 <= '1';
		else
		 s_Energy_Bin_Pos_337 <= s_Energy_Bin_Pos_337;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_337 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_337;   
  
  Energy_Bin_Pos_338 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_338   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_338 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E338_C1_L_Pos and PEAK_C1_Pos <= s_E338_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_338 <= s_Energy_Bin_Pos_338 +'1';
		 Energy_Bin_Pos_Rdy_338 <= '1';
		else
		 s_Energy_Bin_Pos_338 <= s_Energy_Bin_Pos_338;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_338 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_338;   
  
  Energy_Bin_Pos_339 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_339   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_339 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E339_C1_L_Pos and PEAK_C1_Pos <= s_E339_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_339 <= s_Energy_Bin_Pos_339 +'1';
		 Energy_Bin_Pos_Rdy_339 <= '1';
		else
		 s_Energy_Bin_Pos_339 <= s_Energy_Bin_Pos_339;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_339 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_339;         
  
     Energy_Bin_Pos_340 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_340   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_340 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E340_C1_L_Pos and PEAK_C1_Pos <= s_E340_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_340 <= s_Energy_Bin_Pos_340 +'1';
		 Energy_Bin_Pos_Rdy_340 <= '1';
		else
		 s_Energy_Bin_Pos_340 <= s_Energy_Bin_Pos_340;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_340 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_340;    
  
  Energy_Bin_Pos_341 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_341   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_341 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E341_C1_L_Pos and PEAK_C1_Pos <= s_E341_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_341 <= s_Energy_Bin_Pos_341 +'1';
		 Energy_Bin_Pos_Rdy_341 <= '1';
		else
		 s_Energy_Bin_Pos_341 <= s_Energy_Bin_Pos_341;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_341 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_341;   
  
  Energy_Bin_Pos_342 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_342   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_342 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E342_C1_L_Pos and PEAK_C1_Pos <= s_E342_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_342 <= s_Energy_Bin_Pos_342 +'1';
		 Energy_Bin_Pos_Rdy_342 <= '1';
		else
		 s_Energy_Bin_Pos_342 <= s_Energy_Bin_Pos_342;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_342 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_342;   
  
  Energy_Bin_Pos_343 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_343   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_343 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E343_C1_L_Pos and PEAK_C1_Pos <= s_E343_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_343 <= s_Energy_Bin_Pos_343 +'1';
		 Energy_Bin_Pos_Rdy_343 <= '1';
		else
		 s_Energy_Bin_Pos_343 <= s_Energy_Bin_Pos_343;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_343 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_343;   
  
  Energy_Bin_Pos_344 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_344   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_344 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E344_C1_L_Pos and PEAK_C1_Pos <= s_E344_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_344 <= s_Energy_Bin_Pos_344 +'1';
		 Energy_Bin_Pos_Rdy_344 <= '1';
		else
		 s_Energy_Bin_Pos_344 <= s_Energy_Bin_Pos_344;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_344 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_344;   
 
 
  Energy_Bin_Pos_345 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_345   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_345 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E345_C1_L_Pos and PEAK_C1_Pos <= s_E345_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_345 <= s_Energy_Bin_Pos_345 +'1';
		 Energy_Bin_Pos_Rdy_345 <= '1';
		else
		 s_Energy_Bin_Pos_345 <= s_Energy_Bin_Pos_345;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_345 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_345;  
 
  
  Energy_Bin_Pos_346 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_346   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_346 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E346_C1_L_Pos and PEAK_C1_Pos <= s_E346_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_346 <= s_Energy_Bin_Pos_346 +'1';
		 Energy_Bin_Pos_Rdy_346 <= '1';
		else
		 s_Energy_Bin_Pos_346 <= s_Energy_Bin_Pos_346;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_346 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_346;   
  
 Energy_Bin_Pos_347 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_347   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_347 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E347_C1_L_Pos and PEAK_C1_Pos <= s_E347_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_347 <= s_Energy_Bin_Pos_347 +'1';
		 Energy_Bin_Pos_Rdy_347 <= '1';
		else
		 s_Energy_Bin_Pos_347 <= s_Energy_Bin_Pos_347;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_347 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_347;   
  
  Energy_Bin_Pos_348 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_348   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_348 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E348_C1_L_Pos and PEAK_C1_Pos <= s_E348_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_348 <= s_Energy_Bin_Pos_348 +'1';
		 Energy_Bin_Pos_Rdy_348 <= '1';
		else
		 s_Energy_Bin_Pos_348 <= s_Energy_Bin_Pos_348;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_348 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_348;   
  
  Energy_Bin_Pos_349 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_349   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_349 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E349_C1_L_Pos and PEAK_C1_Pos <= s_E349_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_349 <= s_Energy_Bin_Pos_349 +'1';
		 Energy_Bin_Pos_Rdy_349 <= '1';
		else
		 s_Energy_Bin_Pos_349 <= s_Energy_Bin_Pos_349;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_349 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_349;          
  
  
     Energy_Bin_Pos_350 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_350   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_350 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E350_C1_L_Pos and PEAK_C1_Pos <= s_E350_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_350 <= s_Energy_Bin_Pos_350 +'1';
		 Energy_Bin_Pos_Rdy_350 <= '1';
		else
		 s_Energy_Bin_Pos_350 <= s_Energy_Bin_Pos_350;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_350 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_350;    
  
  Energy_Bin_Pos_351 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_351   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_351 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E351_C1_L_Pos and PEAK_C1_Pos <= s_E351_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_351 <= s_Energy_Bin_Pos_351 +'1';
		 Energy_Bin_Pos_Rdy_351 <= '1';
		else
		 s_Energy_Bin_Pos_351 <= s_Energy_Bin_Pos_351;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_351 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_351;   
  
  Energy_Bin_Pos_352 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_352   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_352 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E352_C1_L_Pos and PEAK_C1_Pos <= s_E352_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_352 <= s_Energy_Bin_Pos_352 +'1';
		 Energy_Bin_Pos_Rdy_352 <= '1';
		else
		 s_Energy_Bin_Pos_352 <= s_Energy_Bin_Pos_352;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_352 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_352;   
  
  Energy_Bin_Pos_353 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_353   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_353 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E353_C1_L_Pos and PEAK_C1_Pos <= s_E353_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_353 <= s_Energy_Bin_Pos_353 +'1';
		 Energy_Bin_Pos_Rdy_353 <= '1';
		else
		 s_Energy_Bin_Pos_353 <= s_Energy_Bin_Pos_353;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_353 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_353;   
  
  Energy_Bin_Pos_354 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_354   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_354 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E354_C1_L_Pos and PEAK_C1_Pos <= s_E354_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_354 <= s_Energy_Bin_Pos_354 +'1';
		 Energy_Bin_Pos_Rdy_354 <= '1';
		else
		 s_Energy_Bin_Pos_354 <= s_Energy_Bin_Pos_354;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_354 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_354;   
 
 
  Energy_Bin_Pos_355 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_355   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_355 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E355_C1_L_Pos and PEAK_C1_Pos <= s_E355_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_355 <= s_Energy_Bin_Pos_355 +'1';
		 Energy_Bin_Pos_Rdy_355 <= '1';
		else
		 s_Energy_Bin_Pos_355 <= s_Energy_Bin_Pos_355;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_355 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_355;  
 
  
  Energy_Bin_Pos_356 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_356   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_356 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E356_C1_L_Pos and PEAK_C1_Pos <= s_E356_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_356 <= s_Energy_Bin_Pos_356 +'1';
		 Energy_Bin_Pos_Rdy_356 <= '1';
		else
		 s_Energy_Bin_Pos_356 <= s_Energy_Bin_Pos_356;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_356 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_356;   
  
 Energy_Bin_Pos_357 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_357   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_357 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E357_C1_L_Pos and PEAK_C1_Pos <= s_E357_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_357 <= s_Energy_Bin_Pos_357 +'1';
		 Energy_Bin_Pos_Rdy_357 <= '1';
		else
		 s_Energy_Bin_Pos_357 <= s_Energy_Bin_Pos_357;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_357 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_357;   
  
  Energy_Bin_Pos_358 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_358   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_358 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E358_C1_L_Pos and PEAK_C1_Pos <= s_E358_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_358 <= s_Energy_Bin_Pos_358 +'1';
		 Energy_Bin_Pos_Rdy_358 <= '1';
		else
		 s_Energy_Bin_Pos_358 <= s_Energy_Bin_Pos_358;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_358 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_358;   
  
  Energy_Bin_Pos_359 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_359   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_359 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E359_C1_L_Pos and PEAK_C1_Pos <= s_E359_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_359 <= s_Energy_Bin_Pos_359 +'1';
		 Energy_Bin_Pos_Rdy_359 <= '1';
		else
		 s_Energy_Bin_Pos_359 <= s_Energy_Bin_Pos_359;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_359 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_359;           
  
     Energy_Bin_Pos_360 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_360   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_360 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E360_C1_L_Pos and PEAK_C1_Pos <= s_E360_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_360 <= s_Energy_Bin_Pos_360 +'1';
		 Energy_Bin_Pos_Rdy_360 <= '1';
		else
		 s_Energy_Bin_Pos_360 <= s_Energy_Bin_Pos_360;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_360 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_360;    
  
  Energy_Bin_Pos_361 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_361   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_361 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E361_C1_L_Pos and PEAK_C1_Pos <= s_E361_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_361 <= s_Energy_Bin_Pos_361 +'1';
		 Energy_Bin_Pos_Rdy_361 <= '1';
		else
		 s_Energy_Bin_Pos_361 <= s_Energy_Bin_Pos_361;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_361 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_361;   
  
  Energy_Bin_Pos_362 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_362   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_362 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E362_C1_L_Pos and PEAK_C1_Pos <= s_E362_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_362 <= s_Energy_Bin_Pos_362 +'1';
		 Energy_Bin_Pos_Rdy_362 <= '1';
		else
		 s_Energy_Bin_Pos_362 <= s_Energy_Bin_Pos_362;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_362 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_362;   
  
  Energy_Bin_Pos_363 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_363   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_363 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E363_C1_L_Pos and PEAK_C1_Pos <= s_E363_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_363 <= s_Energy_Bin_Pos_363 +'1';
		 Energy_Bin_Pos_Rdy_363 <= '1';
		else
		 s_Energy_Bin_Pos_363 <= s_Energy_Bin_Pos_363;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_363 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_363;   
  
  Energy_Bin_Pos_364 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_364   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_364 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E364_C1_L_Pos and PEAK_C1_Pos <= s_E364_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_364 <= s_Energy_Bin_Pos_364 +'1';
		 Energy_Bin_Pos_Rdy_364 <= '1';
		else
		 s_Energy_Bin_Pos_364 <= s_Energy_Bin_Pos_364;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_364 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_364;   
 
 
  Energy_Bin_Pos_365 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_365   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_365 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E365_C1_L_Pos and PEAK_C1_Pos <= s_E365_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_365 <= s_Energy_Bin_Pos_365 +'1';
		 Energy_Bin_Pos_Rdy_365 <= '1';
		else
		 s_Energy_Bin_Pos_365 <= s_Energy_Bin_Pos_365;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_365 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_365;  
 
  
  Energy_Bin_Pos_366 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_366   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_366 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E366_C1_L_Pos and PEAK_C1_Pos <= s_E366_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_366 <= s_Energy_Bin_Pos_366 +'1';
		 Energy_Bin_Pos_Rdy_366 <= '1';
		else
		 s_Energy_Bin_Pos_366 <= s_Energy_Bin_Pos_366;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_366 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_366;   
  
 Energy_Bin_Pos_367 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_367   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_367 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E367_C1_L_Pos and PEAK_C1_Pos <= s_E367_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_367 <= s_Energy_Bin_Pos_367 +'1';
		 Energy_Bin_Pos_Rdy_367 <= '1';
		else
		 s_Energy_Bin_Pos_367 <= s_Energy_Bin_Pos_367;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_367 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_367;   
  
  Energy_Bin_Pos_368 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_368   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_368 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E368_C1_L_Pos and PEAK_C1_Pos <= s_E368_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_368 <= s_Energy_Bin_Pos_368 +'1';
		 Energy_Bin_Pos_Rdy_368 <= '1';
		else
		 s_Energy_Bin_Pos_368 <= s_Energy_Bin_Pos_368;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_368 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_368;   
  
  Energy_Bin_Pos_369 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_369   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_369 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E369_C1_L_Pos and PEAK_C1_Pos <= s_E369_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_369 <= s_Energy_Bin_Pos_369 +'1';
		 Energy_Bin_Pos_Rdy_369 <= '1';
		else
		 s_Energy_Bin_Pos_369 <= s_Energy_Bin_Pos_369;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_369 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_369;         
  
     Energy_Bin_Pos_370 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_370   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_370 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E370_C1_L_Pos and PEAK_C1_Pos <= s_E370_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_370 <= s_Energy_Bin_Pos_370 +'1';
		 Energy_Bin_Pos_Rdy_370 <= '1';
		else
		 s_Energy_Bin_Pos_370 <= s_Energy_Bin_Pos_370;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_370 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_370;    
  
  Energy_Bin_Pos_371 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_371   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_371 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E371_C1_L_Pos and PEAK_C1_Pos <= s_E371_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_371 <= s_Energy_Bin_Pos_371 +'1';
		 Energy_Bin_Pos_Rdy_371 <= '1';
		else
		 s_Energy_Bin_Pos_371 <= s_Energy_Bin_Pos_371;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_371 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_371;   
  
  Energy_Bin_Pos_372 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_372   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_372 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E372_C1_L_Pos and PEAK_C1_Pos <= s_E372_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_372 <= s_Energy_Bin_Pos_372 +'1';
		 Energy_Bin_Pos_Rdy_372 <= '1';
		else
		 s_Energy_Bin_Pos_372 <= s_Energy_Bin_Pos_372;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_372 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_372;   
  
  Energy_Bin_Pos_373 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_373   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_373 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E373_C1_L_Pos and PEAK_C1_Pos <= s_E373_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_373 <= s_Energy_Bin_Pos_373 +'1';
		 Energy_Bin_Pos_Rdy_373 <= '1';
		else
		 s_Energy_Bin_Pos_373 <= s_Energy_Bin_Pos_373;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_373 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_373;   
  
  Energy_Bin_Pos_374 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_374   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_374 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E374_C1_L_Pos and PEAK_C1_Pos <= s_E374_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_374 <= s_Energy_Bin_Pos_374 +'1';
		 Energy_Bin_Pos_Rdy_374 <= '1';
		else
		 s_Energy_Bin_Pos_374 <= s_Energy_Bin_Pos_374;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_374 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_374;   
 
 
  Energy_Bin_Pos_375 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_375   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_375 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E375_C1_L_Pos and PEAK_C1_Pos <= s_E375_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_375 <= s_Energy_Bin_Pos_375 +'1';
		 Energy_Bin_Pos_Rdy_375 <= '1';
		else
		 s_Energy_Bin_Pos_375 <= s_Energy_Bin_Pos_375;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_375 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_375;  
 
  
  Energy_Bin_Pos_376 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_376   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_376 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E376_C1_L_Pos and PEAK_C1_Pos <= s_E376_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_376 <= s_Energy_Bin_Pos_376 +'1';
		 Energy_Bin_Pos_Rdy_376 <= '1';
		else
		 s_Energy_Bin_Pos_376 <= s_Energy_Bin_Pos_376;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_376 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_376;   
  
 Energy_Bin_Pos_377 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_377   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_377 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E377_C1_L_Pos and PEAK_C1_Pos <= s_E377_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_377 <= s_Energy_Bin_Pos_377 +'1';
		 Energy_Bin_Pos_Rdy_377 <= '1';
		else
		 s_Energy_Bin_Pos_377 <= s_Energy_Bin_Pos_377;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_377 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_377;   
  
  Energy_Bin_Pos_378 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_378   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_378 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E378_C1_L_Pos and PEAK_C1_Pos <= s_E378_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_378 <= s_Energy_Bin_Pos_378 +'1';
		 Energy_Bin_Pos_Rdy_378 <= '1';
		else
		 s_Energy_Bin_Pos_378 <= s_Energy_Bin_Pos_378;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_378 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_378;   
  
  Energy_Bin_Pos_379 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_379   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_379 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E379_C1_L_Pos and PEAK_C1_Pos <= s_E379_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_379 <= s_Energy_Bin_Pos_379 +'1';
		 Energy_Bin_Pos_Rdy_379 <= '1';
		else
		 s_Energy_Bin_Pos_379 <= s_Energy_Bin_Pos_379;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_379 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_379;       
  
     Energy_Bin_Pos_380 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_380   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_380 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E380_C1_L_Pos and PEAK_C1_Pos <= s_E380_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_380 <= s_Energy_Bin_Pos_380 +'1';
		 Energy_Bin_Pos_Rdy_380 <= '1';
		else
		 s_Energy_Bin_Pos_380 <= s_Energy_Bin_Pos_380;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_380 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_380;    
  
  Energy_Bin_Pos_381 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_381   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_381 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E381_C1_L_Pos and PEAK_C1_Pos <= s_E381_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_381 <= s_Energy_Bin_Pos_381 +'1';
		 Energy_Bin_Pos_Rdy_381 <= '1';
		else
		 s_Energy_Bin_Pos_381 <= s_Energy_Bin_Pos_381;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_381 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_381;   
  
  Energy_Bin_Pos_382 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_382   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_382 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E382_C1_L_Pos and PEAK_C1_Pos <= s_E382_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_382 <= s_Energy_Bin_Pos_382 +'1';
		 Energy_Bin_Pos_Rdy_382 <= '1';
		else
		 s_Energy_Bin_Pos_382 <= s_Energy_Bin_Pos_382;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_382 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_382;   
  
  Energy_Bin_Pos_383 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_383   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_383 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E383_C1_L_Pos and PEAK_C1_Pos <= s_E383_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_383 <= s_Energy_Bin_Pos_383 +'1';
		 Energy_Bin_Pos_Rdy_383 <= '1';
		else
		 s_Energy_Bin_Pos_383 <= s_Energy_Bin_Pos_383;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_383 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_383;   
  
  Energy_Bin_Pos_384 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_384   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_384 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E384_C1_L_Pos and PEAK_C1_Pos <= s_E384_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_384 <= s_Energy_Bin_Pos_384 +'1';
		 Energy_Bin_Pos_Rdy_384 <= '1';
		else
		 s_Energy_Bin_Pos_384 <= s_Energy_Bin_Pos_384;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_384 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_384;   
 
 
  Energy_Bin_Pos_385 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_385   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_385 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E385_C1_L_Pos and PEAK_C1_Pos <= s_E385_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_385 <= s_Energy_Bin_Pos_385 +'1';
		 Energy_Bin_Pos_Rdy_385 <= '1';
		else
		 s_Energy_Bin_Pos_385 <= s_Energy_Bin_Pos_385;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_385 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_385;  
 
  
  Energy_Bin_Pos_386 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_386   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_386 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E386_C1_L_Pos and PEAK_C1_Pos <= s_E386_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_386 <= s_Energy_Bin_Pos_386 +'1';
		 Energy_Bin_Pos_Rdy_386 <= '1';
		else
		 s_Energy_Bin_Pos_386 <= s_Energy_Bin_Pos_386;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_386 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_386;   
  
 Energy_Bin_Pos_387 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_387   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_387 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E387_C1_L_Pos and PEAK_C1_Pos <= s_E387_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_387 <= s_Energy_Bin_Pos_387 +'1';
		 Energy_Bin_Pos_Rdy_387 <= '1';
		else
		 s_Energy_Bin_Pos_387 <= s_Energy_Bin_Pos_387;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_387 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_387;   
  
  Energy_Bin_Pos_388 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_388   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_388 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E388_C1_L_Pos and PEAK_C1_Pos <= s_E388_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_388 <= s_Energy_Bin_Pos_388 +'1';
		 Energy_Bin_Pos_Rdy_388 <= '1';
		else
		 s_Energy_Bin_Pos_388 <= s_Energy_Bin_Pos_388;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_388 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_388;   
  
  Energy_Bin_Pos_389 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_389   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_389 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E389_C1_L_Pos and PEAK_C1_Pos <= s_E389_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_389 <= s_Energy_Bin_Pos_389 +'1';
		 Energy_Bin_Pos_Rdy_389 <= '1';
		else
		 s_Energy_Bin_Pos_389 <= s_Energy_Bin_Pos_389;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_389 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_389;      
  
     Energy_Bin_Pos_390 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_390   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_390 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E390_C1_L_Pos and PEAK_C1_Pos <= s_E390_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_390 <= s_Energy_Bin_Pos_390 +'1';
		 Energy_Bin_Pos_Rdy_390 <= '1';
		else
		 s_Energy_Bin_Pos_390 <= s_Energy_Bin_Pos_390;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_390 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_390;    
  
  Energy_Bin_Pos_391 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_391   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_391 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E391_C1_L_Pos and PEAK_C1_Pos <= s_E391_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_391 <= s_Energy_Bin_Pos_391 +'1';
		 Energy_Bin_Pos_Rdy_391 <= '1';
		else
		 s_Energy_Bin_Pos_391 <= s_Energy_Bin_Pos_391;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_391 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_391;   
  
  Energy_Bin_Pos_392 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_392   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_392 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E392_C1_L_Pos and PEAK_C1_Pos <= s_E392_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_392 <= s_Energy_Bin_Pos_392 +'1';
		 Energy_Bin_Pos_Rdy_392 <= '1';
		else
		 s_Energy_Bin_Pos_392 <= s_Energy_Bin_Pos_392;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_392 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_392;   
  
  Energy_Bin_Pos_393 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_393   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_393 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E393_C1_L_Pos and PEAK_C1_Pos <= s_E393_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_393 <= s_Energy_Bin_Pos_393 +'1';
		 Energy_Bin_Pos_Rdy_393 <= '1';
		else
		 s_Energy_Bin_Pos_393 <= s_Energy_Bin_Pos_393;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_393 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_393;   
  
  Energy_Bin_Pos_394 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_394   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_394 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E394_C1_L_Pos and PEAK_C1_Pos <= s_E394_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_394 <= s_Energy_Bin_Pos_394 +'1';
		 Energy_Bin_Pos_Rdy_394 <= '1';
		else
		 s_Energy_Bin_Pos_394 <= s_Energy_Bin_Pos_394;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_394 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_394;   
 
 
  Energy_Bin_Pos_395 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_395   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_395 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E395_C1_L_Pos and PEAK_C1_Pos <= s_E395_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_395 <= s_Energy_Bin_Pos_395 +'1';
		 Energy_Bin_Pos_Rdy_395 <= '1';
		else
		 s_Energy_Bin_Pos_395 <= s_Energy_Bin_Pos_395;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_395 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_395;  
 
  
  Energy_Bin_Pos_396 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_396   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_396 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E396_C1_L_Pos and PEAK_C1_Pos <= s_E396_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_396 <= s_Energy_Bin_Pos_396 +'1';
		 Energy_Bin_Pos_Rdy_396 <= '1';
		else
		 s_Energy_Bin_Pos_396 <= s_Energy_Bin_Pos_396;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_396 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_396;   
  
 Energy_Bin_Pos_397 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_397   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_397 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E397_C1_L_Pos and PEAK_C1_Pos <= s_E397_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_397 <= s_Energy_Bin_Pos_397 +'1';
		 Energy_Bin_Pos_Rdy_397 <= '1';
		else
		 s_Energy_Bin_Pos_397 <= s_Energy_Bin_Pos_397;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_397 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_397;   
  
  Energy_Bin_Pos_398 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_398   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_398 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E398_C1_L_Pos and PEAK_C1_Pos <= s_E398_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_398 <= s_Energy_Bin_Pos_398 +'1';
		 Energy_Bin_Pos_Rdy_398 <= '1';
		else
		 s_Energy_Bin_Pos_398 <= s_Energy_Bin_Pos_398;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_398 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_398;   
  
  Energy_Bin_Pos_399 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_399   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_399 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E399_C1_L_Pos and PEAK_C1_Pos <= s_E399_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_399 <= s_Energy_Bin_Pos_399 +'1';
		 Energy_Bin_Pos_Rdy_399 <= '1';
		else
		 s_Energy_Bin_Pos_399 <= s_Energy_Bin_Pos_399;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_399 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_399;      

    Energy_Bin_Pos_400 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_400   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_400 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E400_C1_L_Pos and PEAK_C1_Pos <= s_E400_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_400 <= s_Energy_Bin_Pos_400 +'1';
		 Energy_Bin_Pos_Rdy_400 <= '1';
		else
		 s_Energy_Bin_Pos_400 <= s_Energy_Bin_Pos_400;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_400 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_400;    
  
  Energy_Bin_Pos_401 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_401   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_401 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E401_C1_L_Pos and PEAK_C1_Pos <= s_E401_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_401 <= s_Energy_Bin_Pos_401 +'1';
		 Energy_Bin_Pos_Rdy_401 <= '1';
		else
		 s_Energy_Bin_Pos_401 <= s_Energy_Bin_Pos_401;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_401 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_401;   
  
  Energy_Bin_Pos_402 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_402   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_402 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E402_C1_L_Pos and PEAK_C1_Pos <= s_E402_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_402 <= s_Energy_Bin_Pos_402 +'1';
		 Energy_Bin_Pos_Rdy_402 <= '1';
		else
		 s_Energy_Bin_Pos_402 <= s_Energy_Bin_Pos_402;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_402 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_402;   
  
  Energy_Bin_Pos_403 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_403   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_403 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E403_C1_L_Pos and PEAK_C1_Pos <= s_E403_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_403 <= s_Energy_Bin_Pos_403 +'1';
		 Energy_Bin_Pos_Rdy_403 <= '1';
		else
		 s_Energy_Bin_Pos_403 <= s_Energy_Bin_Pos_403;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_403 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_403;   
  
  Energy_Bin_Pos_404 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_404   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_404 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E404_C1_L_Pos and PEAK_C1_Pos <= s_E404_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_404 <= s_Energy_Bin_Pos_404 +'1';
		 Energy_Bin_Pos_Rdy_404 <= '1';
		else
		 s_Energy_Bin_Pos_404 <= s_Energy_Bin_Pos_404;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_404 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_404;   
 
 
  Energy_Bin_Pos_405 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_405   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_405 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E405_C1_L_Pos and PEAK_C1_Pos <= s_E405_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_405 <= s_Energy_Bin_Pos_405 +'1';
		 Energy_Bin_Pos_Rdy_405 <= '1';
		else
		 s_Energy_Bin_Pos_405 <= s_Energy_Bin_Pos_405;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_405 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_405;  
 
  
  Energy_Bin_Pos_406 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_406   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_406 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E406_C1_L_Pos and PEAK_C1_Pos <= s_E406_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_406 <= s_Energy_Bin_Pos_406 +'1';
		 Energy_Bin_Pos_Rdy_406 <= '1';
		else
		 s_Energy_Bin_Pos_406 <= s_Energy_Bin_Pos_406;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_406 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_406;   
  
 Energy_Bin_Pos_407 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_407   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_407 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E407_C1_L_Pos and PEAK_C1_Pos <= s_E407_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_407 <= s_Energy_Bin_Pos_407 +'1';
		 Energy_Bin_Pos_Rdy_407 <= '1';
		else
		 s_Energy_Bin_Pos_407 <= s_Energy_Bin_Pos_407;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_407 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_407;   
  
  Energy_Bin_Pos_408 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_408   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_408 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E408_C1_L_Pos and PEAK_C1_Pos <= s_E408_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_408 <= s_Energy_Bin_Pos_408 +'1';
		 Energy_Bin_Pos_Rdy_408 <= '1';
		else
		 s_Energy_Bin_Pos_408 <= s_Energy_Bin_Pos_408;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_408 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_408;   
  
  Energy_Bin_Pos_409 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_409   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_409 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E409_C1_L_Pos and PEAK_C1_Pos <= s_E409_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_409 <= s_Energy_Bin_Pos_409 +'1';
		 Energy_Bin_Pos_Rdy_409 <= '1';
		else
		 s_Energy_Bin_Pos_409 <= s_Energy_Bin_Pos_409;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_409 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_409;      
  
     Energy_Bin_Pos_410 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_410   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_410 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E410_C1_L_Pos and PEAK_C1_Pos <= s_E410_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_410 <= s_Energy_Bin_Pos_410 +'1';
		 Energy_Bin_Pos_Rdy_410 <= '1';
		else
		 s_Energy_Bin_Pos_410 <= s_Energy_Bin_Pos_410;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_410 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_410;    
  
  Energy_Bin_Pos_411 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_411   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_411 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E411_C1_L_Pos and PEAK_C1_Pos <= s_E411_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_411 <= s_Energy_Bin_Pos_411 +'1';
		 Energy_Bin_Pos_Rdy_411 <= '1';
		else
		 s_Energy_Bin_Pos_411 <= s_Energy_Bin_Pos_411;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_411 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_411;   
  
  Energy_Bin_Pos_412 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_412   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_412 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E412_C1_L_Pos and PEAK_C1_Pos <= s_E412_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_412 <= s_Energy_Bin_Pos_412 +'1';
		 Energy_Bin_Pos_Rdy_412 <= '1';
		else
		 s_Energy_Bin_Pos_412 <= s_Energy_Bin_Pos_412;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_412 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_412;   
  
  Energy_Bin_Pos_413 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_413   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_413 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E413_C1_L_Pos and PEAK_C1_Pos <= s_E413_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_413 <= s_Energy_Bin_Pos_413 +'1';
		 Energy_Bin_Pos_Rdy_413 <= '1';
		else
		 s_Energy_Bin_Pos_413 <= s_Energy_Bin_Pos_413;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_413 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_413;   
  
  Energy_Bin_Pos_414 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_414   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_414 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E414_C1_L_Pos and PEAK_C1_Pos <= s_E414_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_414 <= s_Energy_Bin_Pos_414 +'1';
		 Energy_Bin_Pos_Rdy_414 <= '1';
		else
		 s_Energy_Bin_Pos_414 <= s_Energy_Bin_Pos_414;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_414 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_414;   
 
 
  Energy_Bin_Pos_415 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_415   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_415 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E415_C1_L_Pos and PEAK_C1_Pos <= s_E415_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_415 <= s_Energy_Bin_Pos_415 +'1';
		 Energy_Bin_Pos_Rdy_415 <= '1';
		else
		 s_Energy_Bin_Pos_415 <= s_Energy_Bin_Pos_415;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_415 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_415;  
 
  
  Energy_Bin_Pos_416 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_416   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_416 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E416_C1_L_Pos and PEAK_C1_Pos <= s_E416_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_416 <= s_Energy_Bin_Pos_416 +'1';
		 Energy_Bin_Pos_Rdy_416 <= '1';
		else
		 s_Energy_Bin_Pos_416 <= s_Energy_Bin_Pos_416;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_416 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_416;   
  
 Energy_Bin_Pos_417 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_417   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_417 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E417_C1_L_Pos and PEAK_C1_Pos <= s_E417_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_417 <= s_Energy_Bin_Pos_417 +'1';
		 Energy_Bin_Pos_Rdy_417 <= '1';
		else
		 s_Energy_Bin_Pos_417 <= s_Energy_Bin_Pos_417;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_417 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_417;   
  
  Energy_Bin_Pos_418 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_418   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_418 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E418_C1_L_Pos and PEAK_C1_Pos <= s_E418_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_418 <= s_Energy_Bin_Pos_418 +'1';
		 Energy_Bin_Pos_Rdy_418 <= '1';
		else
		 s_Energy_Bin_Pos_418 <= s_Energy_Bin_Pos_418;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_418 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_418;   
  
  Energy_Bin_Pos_419 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_419   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_419 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E419_C1_L_Pos and PEAK_C1_Pos <= s_E419_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_419 <= s_Energy_Bin_Pos_419 +'1';
		 Energy_Bin_Pos_Rdy_419 <= '1';
		else
		 s_Energy_Bin_Pos_419 <= s_Energy_Bin_Pos_419;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_419 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_419;       
  
     Energy_Bin_Pos_420 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_420   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_420 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E420_C1_L_Pos and PEAK_C1_Pos <= s_E420_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_420 <= s_Energy_Bin_Pos_420 +'1';
		 Energy_Bin_Pos_Rdy_420 <= '1';
		else
		 s_Energy_Bin_Pos_420 <= s_Energy_Bin_Pos_420;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_420 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_420;    
  
  Energy_Bin_Pos_421 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_421   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_421 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E421_C1_L_Pos and PEAK_C1_Pos <= s_E421_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_421 <= s_Energy_Bin_Pos_421 +'1';
		 Energy_Bin_Pos_Rdy_421 <= '1';
		else
		 s_Energy_Bin_Pos_421 <= s_Energy_Bin_Pos_421;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_421 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_421;   
  
  Energy_Bin_Pos_422 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_422   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_422 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E422_C1_L_Pos and PEAK_C1_Pos <= s_E422_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_422 <= s_Energy_Bin_Pos_422 +'1';
		 Energy_Bin_Pos_Rdy_422 <= '1';
		else
		 s_Energy_Bin_Pos_422 <= s_Energy_Bin_Pos_422;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_422 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_422;   
  
  Energy_Bin_Pos_423 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_423   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_423 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E423_C1_L_Pos and PEAK_C1_Pos <= s_E423_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_423 <= s_Energy_Bin_Pos_423 +'1';
		 Energy_Bin_Pos_Rdy_423 <= '1';
		else
		 s_Energy_Bin_Pos_423 <= s_Energy_Bin_Pos_423;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_423 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_423;   
  
  Energy_Bin_Pos_424 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_424   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_424 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E424_C1_L_Pos and PEAK_C1_Pos <= s_E424_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_424 <= s_Energy_Bin_Pos_424 +'1';
		 Energy_Bin_Pos_Rdy_424 <= '1';
		else
		 s_Energy_Bin_Pos_424 <= s_Energy_Bin_Pos_424;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_424 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_424;   
 
 
  Energy_Bin_Pos_425 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_425   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_425 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E425_C1_L_Pos and PEAK_C1_Pos <= s_E425_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_425 <= s_Energy_Bin_Pos_425 +'1';
		 Energy_Bin_Pos_Rdy_425 <= '1';
		else
		 s_Energy_Bin_Pos_425 <= s_Energy_Bin_Pos_425;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_425 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_425;  
 
  
  Energy_Bin_Pos_426 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_426   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_426 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E426_C1_L_Pos and PEAK_C1_Pos <= s_E426_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_426 <= s_Energy_Bin_Pos_426 +'1';
		 Energy_Bin_Pos_Rdy_426 <= '1';
		else
		 s_Energy_Bin_Pos_426 <= s_Energy_Bin_Pos_426;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_426 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_426;   
  
 Energy_Bin_Pos_427 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_427   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_427 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E427_C1_L_Pos and PEAK_C1_Pos <= s_E427_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_427 <= s_Energy_Bin_Pos_427 +'1';
		 Energy_Bin_Pos_Rdy_427 <= '1';
		else
		 s_Energy_Bin_Pos_427 <= s_Energy_Bin_Pos_427;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_427 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_427;   
  
  Energy_Bin_Pos_428 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_428   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_428 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E428_C1_L_Pos and PEAK_C1_Pos <= s_E428_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_428 <= s_Energy_Bin_Pos_428 +'1';
		 Energy_Bin_Pos_Rdy_428 <= '1';
		else
		 s_Energy_Bin_Pos_428 <= s_Energy_Bin_Pos_428;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_428 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_428;   
  
  Energy_Bin_Pos_429 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_429   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_429 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E429_C1_L_Pos and PEAK_C1_Pos <= s_E429_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_429 <= s_Energy_Bin_Pos_429 +'1';
		 Energy_Bin_Pos_Rdy_429 <= '1';
		else
		 s_Energy_Bin_Pos_429 <= s_Energy_Bin_Pos_429;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_429 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_429;        
  
     Energy_Bin_Pos_430 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_430   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_430 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E430_C1_L_Pos and PEAK_C1_Pos <= s_E430_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_430 <= s_Energy_Bin_Pos_430 +'1';
		 Energy_Bin_Pos_Rdy_430 <= '1';
		else
		 s_Energy_Bin_Pos_430 <= s_Energy_Bin_Pos_430;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_430 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_430;    
  
  Energy_Bin_Pos_431 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_431   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_431 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E431_C1_L_Pos and PEAK_C1_Pos <= s_E431_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_431 <= s_Energy_Bin_Pos_431 +'1';
		 Energy_Bin_Pos_Rdy_431 <= '1';
		else
		 s_Energy_Bin_Pos_431 <= s_Energy_Bin_Pos_431;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_431 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_431;   
  
  Energy_Bin_Pos_432 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_432   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_432 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E432_C1_L_Pos and PEAK_C1_Pos <= s_E432_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_432 <= s_Energy_Bin_Pos_432 +'1';
		 Energy_Bin_Pos_Rdy_432 <= '1';
		else
		 s_Energy_Bin_Pos_432 <= s_Energy_Bin_Pos_432;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_432 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_432;   
  
  Energy_Bin_Pos_433 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_433   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_433 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E433_C1_L_Pos and PEAK_C1_Pos <= s_E433_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_433 <= s_Energy_Bin_Pos_433 +'1';
		 Energy_Bin_Pos_Rdy_433 <= '1';
		else
		 s_Energy_Bin_Pos_433 <= s_Energy_Bin_Pos_433;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_433 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_433;   
  
  Energy_Bin_Pos_434 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_434   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_434 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E434_C1_L_Pos and PEAK_C1_Pos <= s_E434_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_434 <= s_Energy_Bin_Pos_434 +'1';
		 Energy_Bin_Pos_Rdy_434 <= '1';
		else
		 s_Energy_Bin_Pos_434 <= s_Energy_Bin_Pos_434;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_434 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_434;   
 
 
  Energy_Bin_Pos_435 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_435   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_435 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E435_C1_L_Pos and PEAK_C1_Pos <= s_E435_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_435 <= s_Energy_Bin_Pos_435 +'1';
		 Energy_Bin_Pos_Rdy_435 <= '1';
		else
		 s_Energy_Bin_Pos_435 <= s_Energy_Bin_Pos_435;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_435 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_435;  
 
  
  Energy_Bin_Pos_436 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_436   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_436 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E436_C1_L_Pos and PEAK_C1_Pos <= s_E436_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_436 <= s_Energy_Bin_Pos_436 +'1';
		 Energy_Bin_Pos_Rdy_436 <= '1';
		else
		 s_Energy_Bin_Pos_436 <= s_Energy_Bin_Pos_436;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_436 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_436;   
  
 Energy_Bin_Pos_437 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_437   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_437 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E437_C1_L_Pos and PEAK_C1_Pos <= s_E437_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_437 <= s_Energy_Bin_Pos_437 +'1';
		 Energy_Bin_Pos_Rdy_437 <= '1';
		else
		 s_Energy_Bin_Pos_437 <= s_Energy_Bin_Pos_437;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_437 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_437;   
  
  Energy_Bin_Pos_438 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_438   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_438 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E438_C1_L_Pos and PEAK_C1_Pos <= s_E438_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_438 <= s_Energy_Bin_Pos_438 +'1';
		 Energy_Bin_Pos_Rdy_438 <= '1';
		else
		 s_Energy_Bin_Pos_438 <= s_Energy_Bin_Pos_438;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_438 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_438;   
  
  Energy_Bin_Pos_439 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_439   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_439 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E439_C1_L_Pos and PEAK_C1_Pos <= s_E439_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_439 <= s_Energy_Bin_Pos_439 +'1';
		 Energy_Bin_Pos_Rdy_439 <= '1';
		else
		 s_Energy_Bin_Pos_439 <= s_Energy_Bin_Pos_439;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_439 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_439;         
  
     Energy_Bin_Pos_440 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_440   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_440 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E440_C1_L_Pos and PEAK_C1_Pos <= s_E440_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_440 <= s_Energy_Bin_Pos_440 +'1';
		 Energy_Bin_Pos_Rdy_440 <= '1';
		else
		 s_Energy_Bin_Pos_440 <= s_Energy_Bin_Pos_440;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_440 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_440;    
  
  Energy_Bin_Pos_441 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_441   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_441 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E441_C1_L_Pos and PEAK_C1_Pos <= s_E441_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_441 <= s_Energy_Bin_Pos_441 +'1';
		 Energy_Bin_Pos_Rdy_441 <= '1';
		else
		 s_Energy_Bin_Pos_441 <= s_Energy_Bin_Pos_441;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_441 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_441;   
  
  Energy_Bin_Pos_442 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_442   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_442 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E442_C1_L_Pos and PEAK_C1_Pos <= s_E442_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_442 <= s_Energy_Bin_Pos_442 +'1';
		 Energy_Bin_Pos_Rdy_442 <= '1';
		else
		 s_Energy_Bin_Pos_442 <= s_Energy_Bin_Pos_442;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_442 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_442;   
  
  Energy_Bin_Pos_443 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_443   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_443 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E443_C1_L_Pos and PEAK_C1_Pos <= s_E443_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_443 <= s_Energy_Bin_Pos_443 +'1';
		 Energy_Bin_Pos_Rdy_443 <= '1';
		else
		 s_Energy_Bin_Pos_443 <= s_Energy_Bin_Pos_443;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_443 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_443;   
  
  Energy_Bin_Pos_444 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_444   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_444 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E444_C1_L_Pos and PEAK_C1_Pos <= s_E444_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_444 <= s_Energy_Bin_Pos_444 +'1';
		 Energy_Bin_Pos_Rdy_444 <= '1';
		else
		 s_Energy_Bin_Pos_444 <= s_Energy_Bin_Pos_444;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_444 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_444;   
 
 
  Energy_Bin_Pos_445 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_445   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_445 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E445_C1_L_Pos and PEAK_C1_Pos <= s_E445_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_445 <= s_Energy_Bin_Pos_445 +'1';
		 Energy_Bin_Pos_Rdy_445 <= '1';
		else
		 s_Energy_Bin_Pos_445 <= s_Energy_Bin_Pos_445;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_445 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_445;  
 
  
  Energy_Bin_Pos_446 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_446   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_446 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E446_C1_L_Pos and PEAK_C1_Pos <= s_E446_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_446 <= s_Energy_Bin_Pos_446 +'1';
		 Energy_Bin_Pos_Rdy_446 <= '1';
		else
		 s_Energy_Bin_Pos_446 <= s_Energy_Bin_Pos_446;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_446 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_446;   
  
 Energy_Bin_Pos_447 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_447   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_447 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E447_C1_L_Pos and PEAK_C1_Pos <= s_E447_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_447 <= s_Energy_Bin_Pos_447 +'1';
		 Energy_Bin_Pos_Rdy_447 <= '1';
		else
		 s_Energy_Bin_Pos_447 <= s_Energy_Bin_Pos_447;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_447 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_447;   
  
  Energy_Bin_Pos_448 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_448   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_448 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E448_C1_L_Pos and PEAK_C1_Pos <= s_E448_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_448 <= s_Energy_Bin_Pos_448 +'1';
		 Energy_Bin_Pos_Rdy_448 <= '1';
		else
		 s_Energy_Bin_Pos_448 <= s_Energy_Bin_Pos_448;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_448 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_448;   
  
  Energy_Bin_Pos_449 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_449   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_449 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E449_C1_L_Pos and PEAK_C1_Pos <= s_E449_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_449 <= s_Energy_Bin_Pos_449 +'1';
		 Energy_Bin_Pos_Rdy_449 <= '1';
		else
		 s_Energy_Bin_Pos_449 <= s_Energy_Bin_Pos_449;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_449 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_449;          
  
  
     Energy_Bin_Pos_450 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_450   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_450 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E450_C1_L_Pos and PEAK_C1_Pos <= s_E450_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_450 <= s_Energy_Bin_Pos_450 +'1';
		 Energy_Bin_Pos_Rdy_450 <= '1';
		else
		 s_Energy_Bin_Pos_450 <= s_Energy_Bin_Pos_450;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_450 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_450;    
  
  Energy_Bin_Pos_451 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_451   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_451 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E451_C1_L_Pos and PEAK_C1_Pos <= s_E451_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_451 <= s_Energy_Bin_Pos_451 +'1';
		 Energy_Bin_Pos_Rdy_451 <= '1';
		else
		 s_Energy_Bin_Pos_451 <= s_Energy_Bin_Pos_451;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_451 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_451;   
  
  Energy_Bin_Pos_452 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_452   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_452 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E452_C1_L_Pos and PEAK_C1_Pos <= s_E452_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_452 <= s_Energy_Bin_Pos_452 +'1';
		 Energy_Bin_Pos_Rdy_452 <= '1';
		else
		 s_Energy_Bin_Pos_452 <= s_Energy_Bin_Pos_452;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_452 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_452;   
  
  Energy_Bin_Pos_453 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_453   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_453 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E453_C1_L_Pos and PEAK_C1_Pos <= s_E453_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_453 <= s_Energy_Bin_Pos_453 +'1';
		 Energy_Bin_Pos_Rdy_453 <= '1';
		else
		 s_Energy_Bin_Pos_453 <= s_Energy_Bin_Pos_453;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_453 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_453;   
  
  Energy_Bin_Pos_454 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_454   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_454 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E454_C1_L_Pos and PEAK_C1_Pos <= s_E454_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_454 <= s_Energy_Bin_Pos_454 +'1';
		 Energy_Bin_Pos_Rdy_454 <= '1';
		else
		 s_Energy_Bin_Pos_454 <= s_Energy_Bin_Pos_454;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_454 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_454;   
 
 
  Energy_Bin_Pos_455 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_455   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_455 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E455_C1_L_Pos and PEAK_C1_Pos <= s_E455_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_455 <= s_Energy_Bin_Pos_455 +'1';
		 Energy_Bin_Pos_Rdy_455 <= '1';
		else
		 s_Energy_Bin_Pos_455 <= s_Energy_Bin_Pos_455;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_455 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_455;  
 
  
  Energy_Bin_Pos_456 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_456   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_456 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E456_C1_L_Pos and PEAK_C1_Pos <= s_E456_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_456 <= s_Energy_Bin_Pos_456 +'1';
		 Energy_Bin_Pos_Rdy_456 <= '1';
		else
		 s_Energy_Bin_Pos_456 <= s_Energy_Bin_Pos_456;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_456 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_456;   
  
 Energy_Bin_Pos_457 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_457   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_457 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E457_C1_L_Pos and PEAK_C1_Pos <= s_E457_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_457 <= s_Energy_Bin_Pos_457 +'1';
		 Energy_Bin_Pos_Rdy_457 <= '1';
		else
		 s_Energy_Bin_Pos_457 <= s_Energy_Bin_Pos_457;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_457 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_457;   
  
  Energy_Bin_Pos_458 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_458   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_458 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E458_C1_L_Pos and PEAK_C1_Pos <= s_E458_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_458 <= s_Energy_Bin_Pos_458 +'1';
		 Energy_Bin_Pos_Rdy_458 <= '1';
		else
		 s_Energy_Bin_Pos_458 <= s_Energy_Bin_Pos_458;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_458 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_458;   
  
  Energy_Bin_Pos_459 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_459   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_459 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E459_C1_L_Pos and PEAK_C1_Pos <= s_E459_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_459 <= s_Energy_Bin_Pos_459 +'1';
		 Energy_Bin_Pos_Rdy_459 <= '1';
		else
		 s_Energy_Bin_Pos_459 <= s_Energy_Bin_Pos_459;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_459 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_459;           
  
     Energy_Bin_Pos_460 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_460   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_460 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E460_C1_L_Pos and PEAK_C1_Pos <= s_E460_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_460 <= s_Energy_Bin_Pos_460 +'1';
		 Energy_Bin_Pos_Rdy_460 <= '1';
		else
		 s_Energy_Bin_Pos_460 <= s_Energy_Bin_Pos_460;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_460 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_460;    
  
  Energy_Bin_Pos_461 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_461   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_461 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E461_C1_L_Pos and PEAK_C1_Pos <= s_E461_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_461 <= s_Energy_Bin_Pos_461 +'1';
		 Energy_Bin_Pos_Rdy_461 <= '1';
		else
		 s_Energy_Bin_Pos_461 <= s_Energy_Bin_Pos_461;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_461 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_461;   
  
  Energy_Bin_Pos_462 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_462   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_462 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E462_C1_L_Pos and PEAK_C1_Pos <= s_E462_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_462 <= s_Energy_Bin_Pos_462 +'1';
		 Energy_Bin_Pos_Rdy_462 <= '1';
		else
		 s_Energy_Bin_Pos_462 <= s_Energy_Bin_Pos_462;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_462 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_462;   
  
  Energy_Bin_Pos_463 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_463   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_463 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E463_C1_L_Pos and PEAK_C1_Pos <= s_E463_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_463 <= s_Energy_Bin_Pos_463 +'1';
		 Energy_Bin_Pos_Rdy_463 <= '1';
		else
		 s_Energy_Bin_Pos_463 <= s_Energy_Bin_Pos_463;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_463 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_463;   
  
  Energy_Bin_Pos_464 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_464   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_464 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E464_C1_L_Pos and PEAK_C1_Pos <= s_E464_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_464 <= s_Energy_Bin_Pos_464 +'1';
		 Energy_Bin_Pos_Rdy_464 <= '1';
		else
		 s_Energy_Bin_Pos_464 <= s_Energy_Bin_Pos_464;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_464 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_464;   
 
 
  Energy_Bin_Pos_465 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_465   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_465 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E465_C1_L_Pos and PEAK_C1_Pos <= s_E465_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_465 <= s_Energy_Bin_Pos_465 +'1';
		 Energy_Bin_Pos_Rdy_465 <= '1';
		else
		 s_Energy_Bin_Pos_465 <= s_Energy_Bin_Pos_465;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_465 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_465;  
 
  
  Energy_Bin_Pos_466 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_466   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_466 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E466_C1_L_Pos and PEAK_C1_Pos <= s_E466_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_466 <= s_Energy_Bin_Pos_466 +'1';
		 Energy_Bin_Pos_Rdy_466 <= '1';
		else
		 s_Energy_Bin_Pos_466 <= s_Energy_Bin_Pos_466;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_466 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_466;   
  
 Energy_Bin_Pos_467 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_467   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_467 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E467_C1_L_Pos and PEAK_C1_Pos <= s_E467_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_467 <= s_Energy_Bin_Pos_467 +'1';
		 Energy_Bin_Pos_Rdy_467 <= '1';
		else
		 s_Energy_Bin_Pos_467 <= s_Energy_Bin_Pos_467;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_467 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_467;   
  
  Energy_Bin_Pos_468 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_468   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_468 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E468_C1_L_Pos and PEAK_C1_Pos <= s_E468_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_468 <= s_Energy_Bin_Pos_468 +'1';
		 Energy_Bin_Pos_Rdy_468 <= '1';
		else
		 s_Energy_Bin_Pos_468 <= s_Energy_Bin_Pos_468;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_468 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_468;   
  
  Energy_Bin_Pos_469 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_469   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_469 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E469_C1_L_Pos and PEAK_C1_Pos <= s_E469_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_469 <= s_Energy_Bin_Pos_469 +'1';
		 Energy_Bin_Pos_Rdy_469 <= '1';
		else
		 s_Energy_Bin_Pos_469 <= s_Energy_Bin_Pos_469;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_469 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_469;         
  
     Energy_Bin_Pos_470 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_470   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_470 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E470_C1_L_Pos and PEAK_C1_Pos <= s_E470_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_470 <= s_Energy_Bin_Pos_470 +'1';
		 Energy_Bin_Pos_Rdy_470 <= '1';
		else
		 s_Energy_Bin_Pos_470 <= s_Energy_Bin_Pos_470;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_470 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_470;    
  
  Energy_Bin_Pos_471 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_471   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_471 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E471_C1_L_Pos and PEAK_C1_Pos <= s_E471_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_471 <= s_Energy_Bin_Pos_471 +'1';
		 Energy_Bin_Pos_Rdy_471 <= '1';
		else
		 s_Energy_Bin_Pos_471 <= s_Energy_Bin_Pos_471;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_471 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_471;   
  
  Energy_Bin_Pos_472 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_472   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_472 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E472_C1_L_Pos and PEAK_C1_Pos <= s_E472_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_472 <= s_Energy_Bin_Pos_472 +'1';
		 Energy_Bin_Pos_Rdy_472 <= '1';
		else
		 s_Energy_Bin_Pos_472 <= s_Energy_Bin_Pos_472;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_472 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_472;   
  
  Energy_Bin_Pos_473 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_473   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_473 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E473_C1_L_Pos and PEAK_C1_Pos <= s_E473_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_473 <= s_Energy_Bin_Pos_473 +'1';
		 Energy_Bin_Pos_Rdy_473 <= '1';
		else
		 s_Energy_Bin_Pos_473 <= s_Energy_Bin_Pos_473;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_473 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_473;   
  
  Energy_Bin_Pos_474 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_474   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_474 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E474_C1_L_Pos and PEAK_C1_Pos <= s_E474_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_474 <= s_Energy_Bin_Pos_474 +'1';
		 Energy_Bin_Pos_Rdy_474 <= '1';
		else
		 s_Energy_Bin_Pos_474 <= s_Energy_Bin_Pos_474;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_474 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_474;   
 
 
  Energy_Bin_Pos_475 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_475   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_475 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E475_C1_L_Pos and PEAK_C1_Pos <= s_E475_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_475 <= s_Energy_Bin_Pos_475 +'1';
		 Energy_Bin_Pos_Rdy_475 <= '1';
		else
		 s_Energy_Bin_Pos_475 <= s_Energy_Bin_Pos_475;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_475 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_475;  
 
  
  Energy_Bin_Pos_476 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_476   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_476 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E476_C1_L_Pos and PEAK_C1_Pos <= s_E476_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_476 <= s_Energy_Bin_Pos_476 +'1';
		 Energy_Bin_Pos_Rdy_476 <= '1';
		else
		 s_Energy_Bin_Pos_476 <= s_Energy_Bin_Pos_476;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_476 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_476;   
  
 Energy_Bin_Pos_477 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_477   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_477 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E477_C1_L_Pos and PEAK_C1_Pos <= s_E477_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_477 <= s_Energy_Bin_Pos_477 +'1';
		 Energy_Bin_Pos_Rdy_477 <= '1';
		else
		 s_Energy_Bin_Pos_477 <= s_Energy_Bin_Pos_477;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_477 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_477;   
  
  Energy_Bin_Pos_478 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_478   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_478 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E478_C1_L_Pos and PEAK_C1_Pos <= s_E478_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_478 <= s_Energy_Bin_Pos_478 +'1';
		 Energy_Bin_Pos_Rdy_478 <= '1';
		else
		 s_Energy_Bin_Pos_478 <= s_Energy_Bin_Pos_478;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_478 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_478;   
  
  Energy_Bin_Pos_479 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_479   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_479 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E479_C1_L_Pos and PEAK_C1_Pos <= s_E479_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_479 <= s_Energy_Bin_Pos_479 +'1';
		 Energy_Bin_Pos_Rdy_479 <= '1';
		else
		 s_Energy_Bin_Pos_479 <= s_Energy_Bin_Pos_479;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_479 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_479;       
  
     Energy_Bin_Pos_480 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_480   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_480 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E480_C1_L_Pos and PEAK_C1_Pos <= s_E480_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_480 <= s_Energy_Bin_Pos_480 +'1';
		 Energy_Bin_Pos_Rdy_480 <= '1';
		else
		 s_Energy_Bin_Pos_480 <= s_Energy_Bin_Pos_480;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_480 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_480;    
  
  Energy_Bin_Pos_481 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_481   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_481 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E481_C1_L_Pos and PEAK_C1_Pos <= s_E481_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_481 <= s_Energy_Bin_Pos_481 +'1';
		 Energy_Bin_Pos_Rdy_481 <= '1';
		else
		 s_Energy_Bin_Pos_481 <= s_Energy_Bin_Pos_481;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_481 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_481;   
  
  Energy_Bin_Pos_482 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_482   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_482 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E482_C1_L_Pos and PEAK_C1_Pos <= s_E482_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_482 <= s_Energy_Bin_Pos_482 +'1';
		 Energy_Bin_Pos_Rdy_482 <= '1';
		else
		 s_Energy_Bin_Pos_482 <= s_Energy_Bin_Pos_482;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_482 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_482;   
  
  Energy_Bin_Pos_483 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_483   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_483 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E483_C1_L_Pos and PEAK_C1_Pos <= s_E483_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_483 <= s_Energy_Bin_Pos_483 +'1';
		 Energy_Bin_Pos_Rdy_483 <= '1';
		else
		 s_Energy_Bin_Pos_483 <= s_Energy_Bin_Pos_483;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_483 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_483;   
  
  Energy_Bin_Pos_484 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_484   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_484 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E484_C1_L_Pos and PEAK_C1_Pos <= s_E484_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_484 <= s_Energy_Bin_Pos_484 +'1';
		 Energy_Bin_Pos_Rdy_484 <= '1';
		else
		 s_Energy_Bin_Pos_484 <= s_Energy_Bin_Pos_484;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_484 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_484;   
 
 
  Energy_Bin_Pos_485 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_485   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_485 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E485_C1_L_Pos and PEAK_C1_Pos <= s_E485_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_485 <= s_Energy_Bin_Pos_485 +'1';
		 Energy_Bin_Pos_Rdy_485 <= '1';
		else
		 s_Energy_Bin_Pos_485 <= s_Energy_Bin_Pos_485;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_485 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_485;  
 
  
  Energy_Bin_Pos_486 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_486   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_486 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E486_C1_L_Pos and PEAK_C1_Pos <= s_E486_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_486 <= s_Energy_Bin_Pos_486 +'1';
		 Energy_Bin_Pos_Rdy_486 <= '1';
		else
		 s_Energy_Bin_Pos_486 <= s_Energy_Bin_Pos_486;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_486 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_486;   
  
 Energy_Bin_Pos_487 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_487   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_487 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E487_C1_L_Pos and PEAK_C1_Pos <= s_E487_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_487 <= s_Energy_Bin_Pos_487 +'1';
		 Energy_Bin_Pos_Rdy_487 <= '1';
		else
		 s_Energy_Bin_Pos_487 <= s_Energy_Bin_Pos_487;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_487 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_487;   
  
  Energy_Bin_Pos_488 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_488   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_488 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E488_C1_L_Pos and PEAK_C1_Pos <= s_E488_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_488 <= s_Energy_Bin_Pos_488 +'1';
		 Energy_Bin_Pos_Rdy_488 <= '1';
		else
		 s_Energy_Bin_Pos_488 <= s_Energy_Bin_Pos_488;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_488 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_488;   
  
  Energy_Bin_Pos_489 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_489   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_489 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E489_C1_L_Pos and PEAK_C1_Pos <= s_E489_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_489 <= s_Energy_Bin_Pos_489 +'1';
		 Energy_Bin_Pos_Rdy_489 <= '1';
		else
		 s_Energy_Bin_Pos_489 <= s_Energy_Bin_Pos_489;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_489 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_489;      
  
     Energy_Bin_Pos_490 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_490   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_490 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E490_C1_L_Pos and PEAK_C1_Pos <= s_E490_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_490 <= s_Energy_Bin_Pos_490 +'1';
		 Energy_Bin_Pos_Rdy_490 <= '1';
		else
		 s_Energy_Bin_Pos_490 <= s_Energy_Bin_Pos_490;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_490 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_490;    
  
  Energy_Bin_Pos_491 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_491   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_491 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E491_C1_L_Pos and PEAK_C1_Pos <= s_E491_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_491 <= s_Energy_Bin_Pos_491 +'1';
		 Energy_Bin_Pos_Rdy_491 <= '1';
		else
		 s_Energy_Bin_Pos_491 <= s_Energy_Bin_Pos_491;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_491 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_491;   
  
  Energy_Bin_Pos_492 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_492   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_492 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E492_C1_L_Pos and PEAK_C1_Pos <= s_E492_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_492 <= s_Energy_Bin_Pos_492 +'1';
		 Energy_Bin_Pos_Rdy_492 <= '1';
		else
		 s_Energy_Bin_Pos_492 <= s_Energy_Bin_Pos_492;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_492 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_492;   
  
  Energy_Bin_Pos_493 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_493   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_493 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E493_C1_L_Pos and PEAK_C1_Pos <= s_E493_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_493 <= s_Energy_Bin_Pos_493 +'1';
		 Energy_Bin_Pos_Rdy_493 <= '1';
		else
		 s_Energy_Bin_Pos_493 <= s_Energy_Bin_Pos_493;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_493 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_493;   
  
  Energy_Bin_Pos_494 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_494   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_494 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E494_C1_L_Pos and PEAK_C1_Pos <= s_E494_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_494 <= s_Energy_Bin_Pos_494 +'1';
		 Energy_Bin_Pos_Rdy_494 <= '1';
		else
		 s_Energy_Bin_Pos_494 <= s_Energy_Bin_Pos_494;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_494 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_494;   
 
 
  Energy_Bin_Pos_495 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_495   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_495 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E495_C1_L_Pos and PEAK_C1_Pos <= s_E495_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_495 <= s_Energy_Bin_Pos_495 +'1';
		 Energy_Bin_Pos_Rdy_495 <= '1';
		else
		 s_Energy_Bin_Pos_495 <= s_Energy_Bin_Pos_495;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_495 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_495;  
 
  
  Energy_Bin_Pos_496 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_496   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_496 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E496_C1_L_Pos and PEAK_C1_Pos <= s_E496_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_496 <= s_Energy_Bin_Pos_496 +'1';
		 Energy_Bin_Pos_Rdy_496 <= '1';
		else
		 s_Energy_Bin_Pos_496 <= s_Energy_Bin_Pos_496;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_496 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_496;   
  
 Energy_Bin_Pos_497 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_497   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_497 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E497_C1_L_Pos and PEAK_C1_Pos <= s_E497_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_497 <= s_Energy_Bin_Pos_497 +'1';
		 Energy_Bin_Pos_Rdy_497 <= '1';
		else
		 s_Energy_Bin_Pos_497 <= s_Energy_Bin_Pos_497;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_497 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_497;   
  
  Energy_Bin_Pos_498 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_498   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_498 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E498_C1_L_Pos and PEAK_C1_Pos <= s_E498_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_498 <= s_Energy_Bin_Pos_498 +'1';
		 Energy_Bin_Pos_Rdy_498 <= '1';
		else
		 s_Energy_Bin_Pos_498 <= s_Energy_Bin_Pos_498;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_498 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_498;   
  
  Energy_Bin_Pos_499 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_499   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_499 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E499_C1_L_Pos and PEAK_C1_Pos <= s_E499_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_499 <= s_Energy_Bin_Pos_499 +'1';
		 Energy_Bin_Pos_Rdy_499 <= '1';
		else
		 s_Energy_Bin_Pos_499 <= s_Energy_Bin_Pos_499;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_499 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_499;      

    Energy_Bin_Pos_500 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_500   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_500 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E500_C1_L_Pos and PEAK_C1_Pos <= s_E500_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_500 <= s_Energy_Bin_Pos_500 +'1';
		 Energy_Bin_Pos_Rdy_500 <= '1';
		else
		 s_Energy_Bin_Pos_500 <= s_Energy_Bin_Pos_500;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_500 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_500;    
  
  Energy_Bin_Pos_501 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_501   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_501 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E501_C1_L_Pos and PEAK_C1_Pos <= s_E501_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_501 <= s_Energy_Bin_Pos_501 +'1';
		 Energy_Bin_Pos_Rdy_501 <= '1';
		else
		 s_Energy_Bin_Pos_501 <= s_Energy_Bin_Pos_501;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_501 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_501;   
  
  Energy_Bin_Pos_502 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_502   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_502 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E502_C1_L_Pos and PEAK_C1_Pos <= s_E502_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_502 <= s_Energy_Bin_Pos_502 +'1';
		 Energy_Bin_Pos_Rdy_502 <= '1';
		else
		 s_Energy_Bin_Pos_502 <= s_Energy_Bin_Pos_502;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_502 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_502;   
  
  Energy_Bin_Pos_503 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_503   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_503 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E503_C1_L_Pos and PEAK_C1_Pos <= s_E503_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_503 <= s_Energy_Bin_Pos_503 +'1';
		 Energy_Bin_Pos_Rdy_503 <= '1';
		else
		 s_Energy_Bin_Pos_503 <= s_Energy_Bin_Pos_503;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_503 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_503;   
  
  Energy_Bin_Pos_504 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_504   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_504 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E504_C1_L_Pos and PEAK_C1_Pos <= s_E504_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_504 <= s_Energy_Bin_Pos_504 +'1';
		 Energy_Bin_Pos_Rdy_504 <= '1';
		else
		 s_Energy_Bin_Pos_504 <= s_Energy_Bin_Pos_504;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_504 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_504;   
 
 
  Energy_Bin_Pos_505 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_505   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_505 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E505_C1_L_Pos and PEAK_C1_Pos <= s_E505_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_505 <= s_Energy_Bin_Pos_505 +'1';
		 Energy_Bin_Pos_Rdy_505 <= '1';
		else
		 s_Energy_Bin_Pos_505 <= s_Energy_Bin_Pos_505;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_505 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_505;  
 
  
  Energy_Bin_Pos_506 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_506   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_506 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E506_C1_L_Pos and PEAK_C1_Pos <= s_E506_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_506 <= s_Energy_Bin_Pos_506 +'1';
		 Energy_Bin_Pos_Rdy_506 <= '1';
		else
		 s_Energy_Bin_Pos_506 <= s_Energy_Bin_Pos_506;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_506 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_506;   
  
 Energy_Bin_Pos_507 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_507   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_507 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E507_C1_L_Pos and PEAK_C1_Pos <= s_E507_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_507 <= s_Energy_Bin_Pos_507 +'1';
		 Energy_Bin_Pos_Rdy_507 <= '1';
		else
		 s_Energy_Bin_Pos_507 <= s_Energy_Bin_Pos_507;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_507 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_507;   
  
  Energy_Bin_Pos_508 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_508   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_508 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E508_C1_L_Pos and PEAK_C1_Pos <= s_E508_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_508 <= s_Energy_Bin_Pos_508 +'1';
		 Energy_Bin_Pos_Rdy_508 <= '1';
		else
		 s_Energy_Bin_Pos_508 <= s_Energy_Bin_Pos_508;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_508 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_508;   
  
  Energy_Bin_Pos_509 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_509   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_509 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E509_C1_L_Pos and PEAK_C1_Pos <= s_E509_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_509 <= s_Energy_Bin_Pos_509 +'1';
		 Energy_Bin_Pos_Rdy_509 <= '1';
		else
		 s_Energy_Bin_Pos_509 <= s_Energy_Bin_Pos_509;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_509 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_509;      
  
     Energy_Bin_Pos_510 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_510   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_510 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E510_C1_L_Pos and PEAK_C1_Pos <= s_E510_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_510 <= s_Energy_Bin_Pos_510 +'1';
		 Energy_Bin_Pos_Rdy_510 <= '1';
		else
		 s_Energy_Bin_Pos_510 <= s_Energy_Bin_Pos_510;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_510 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_510;    
  
  Energy_Bin_Pos_511 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_511   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_511 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E511_C1_L_Pos and PEAK_C1_Pos <= s_E511_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_511 <= s_Energy_Bin_Pos_511 +'1';
		 Energy_Bin_Pos_Rdy_511 <= '1';
		else
		 s_Energy_Bin_Pos_511 <= s_Energy_Bin_Pos_511;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_511 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_511;   
  
  Energy_Bin_Pos_512 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_512   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_512 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E512_C1_L_Pos and PEAK_C1_Pos <= s_E512_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_512 <= s_Energy_Bin_Pos_512 +'1';
		 Energy_Bin_Pos_Rdy_512 <= '1';
		else
		 s_Energy_Bin_Pos_512 <= s_Energy_Bin_Pos_512;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_512 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_512;   
  
  Energy_Bin_Pos_513 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_513   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_513 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E513_C1_L_Pos and PEAK_C1_Pos <= s_E513_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_513 <= s_Energy_Bin_Pos_513 +'1';
		 Energy_Bin_Pos_Rdy_513 <= '1';
		else
		 s_Energy_Bin_Pos_513 <= s_Energy_Bin_Pos_513;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_513 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_513;   
  
  Energy_Bin_Pos_514 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_514   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_514 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E514_C1_L_Pos and PEAK_C1_Pos <= s_E514_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_514 <= s_Energy_Bin_Pos_514 +'1';
		 Energy_Bin_Pos_Rdy_514 <= '1';
		else
		 s_Energy_Bin_Pos_514 <= s_Energy_Bin_Pos_514;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_514 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_514;   
 
 
  Energy_Bin_Pos_515 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_515   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_515 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E515_C1_L_Pos and PEAK_C1_Pos <= s_E515_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_515 <= s_Energy_Bin_Pos_515 +'1';
		 Energy_Bin_Pos_Rdy_515 <= '1';
		else
		 s_Energy_Bin_Pos_515 <= s_Energy_Bin_Pos_515;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_515 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_515;  
 
  
  Energy_Bin_Pos_516 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_516   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_516 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E516_C1_L_Pos and PEAK_C1_Pos <= s_E516_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_516 <= s_Energy_Bin_Pos_516 +'1';
		 Energy_Bin_Pos_Rdy_516 <= '1';
		else
		 s_Energy_Bin_Pos_516 <= s_Energy_Bin_Pos_516;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_516 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_516;   
  
 Energy_Bin_Pos_517 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_517   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_517 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E517_C1_L_Pos and PEAK_C1_Pos <= s_E517_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_517 <= s_Energy_Bin_Pos_517 +'1';
		 Energy_Bin_Pos_Rdy_517 <= '1';
		else
		 s_Energy_Bin_Pos_517 <= s_Energy_Bin_Pos_517;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_517 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_517;   
  
  Energy_Bin_Pos_518 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_518   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_518 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E518_C1_L_Pos and PEAK_C1_Pos <= s_E518_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_518 <= s_Energy_Bin_Pos_518 +'1';
		 Energy_Bin_Pos_Rdy_518 <= '1';
		else
		 s_Energy_Bin_Pos_518 <= s_Energy_Bin_Pos_518;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_518 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_518;   
  
  Energy_Bin_Pos_519 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_519   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_519 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E519_C1_L_Pos and PEAK_C1_Pos <= s_E519_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_519 <= s_Energy_Bin_Pos_519 +'1';
		 Energy_Bin_Pos_Rdy_519 <= '1';
		else
		 s_Energy_Bin_Pos_519 <= s_Energy_Bin_Pos_519;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_519 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_519;       
  
     Energy_Bin_Pos_520 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_520   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_520 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E520_C1_L_Pos and PEAK_C1_Pos <= s_E520_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_520 <= s_Energy_Bin_Pos_520 +'1';
		 Energy_Bin_Pos_Rdy_520 <= '1';
		else
		 s_Energy_Bin_Pos_520 <= s_Energy_Bin_Pos_520;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_520 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_520;    
  
  Energy_Bin_Pos_521 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_521   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_521 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E521_C1_L_Pos and PEAK_C1_Pos <= s_E521_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_521 <= s_Energy_Bin_Pos_521 +'1';
		 Energy_Bin_Pos_Rdy_521 <= '1';
		else
		 s_Energy_Bin_Pos_521 <= s_Energy_Bin_Pos_521;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_521 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_521;   
  
  Energy_Bin_Pos_522 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_522   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_522 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E522_C1_L_Pos and PEAK_C1_Pos <= s_E522_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_522 <= s_Energy_Bin_Pos_522 +'1';
		 Energy_Bin_Pos_Rdy_522 <= '1';
		else
		 s_Energy_Bin_Pos_522 <= s_Energy_Bin_Pos_522;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_522 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_522;   
  
  Energy_Bin_Pos_523 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_523   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_523 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E523_C1_L_Pos and PEAK_C1_Pos <= s_E523_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_523 <= s_Energy_Bin_Pos_523 +'1';
		 Energy_Bin_Pos_Rdy_523 <= '1';
		else
		 s_Energy_Bin_Pos_523 <= s_Energy_Bin_Pos_523;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_523 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_523;   
  
  Energy_Bin_Pos_524 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_524   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_524 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E524_C1_L_Pos and PEAK_C1_Pos <= s_E524_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_524 <= s_Energy_Bin_Pos_524 +'1';
		 Energy_Bin_Pos_Rdy_524 <= '1';
		else
		 s_Energy_Bin_Pos_524 <= s_Energy_Bin_Pos_524;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_524 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_524;   
 
 
  Energy_Bin_Pos_525 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_525   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_525 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E525_C1_L_Pos and PEAK_C1_Pos <= s_E525_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_525 <= s_Energy_Bin_Pos_525 +'1';
		 Energy_Bin_Pos_Rdy_525 <= '1';
		else
		 s_Energy_Bin_Pos_525 <= s_Energy_Bin_Pos_525;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_525 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_525;  
 
  
  Energy_Bin_Pos_526 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_526   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_526 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E526_C1_L_Pos and PEAK_C1_Pos <= s_E526_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_526 <= s_Energy_Bin_Pos_526 +'1';
		 Energy_Bin_Pos_Rdy_526 <= '1';
		else
		 s_Energy_Bin_Pos_526 <= s_Energy_Bin_Pos_526;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_526 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_526;   
  
 Energy_Bin_Pos_527 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_527   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_527 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E527_C1_L_Pos and PEAK_C1_Pos <= s_E527_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_527 <= s_Energy_Bin_Pos_527 +'1';
		 Energy_Bin_Pos_Rdy_527 <= '1';
		else
		 s_Energy_Bin_Pos_527 <= s_Energy_Bin_Pos_527;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_527 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_527;   
  
  Energy_Bin_Pos_528 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_528   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_528 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E528_C1_L_Pos and PEAK_C1_Pos <= s_E528_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_528 <= s_Energy_Bin_Pos_528 +'1';
		 Energy_Bin_Pos_Rdy_528 <= '1';
		else
		 s_Energy_Bin_Pos_528 <= s_Energy_Bin_Pos_528;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_528 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_528;   
  
  Energy_Bin_Pos_529 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_529   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_529 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E529_C1_L_Pos and PEAK_C1_Pos <= s_E529_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_529 <= s_Energy_Bin_Pos_529 +'1';
		 Energy_Bin_Pos_Rdy_529 <= '1';
		else
		 s_Energy_Bin_Pos_529 <= s_Energy_Bin_Pos_529;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_529 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_529;        
  
     Energy_Bin_Pos_530 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_530   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_530 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E530_C1_L_Pos and PEAK_C1_Pos <= s_E530_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_530 <= s_Energy_Bin_Pos_530 +'1';
		 Energy_Bin_Pos_Rdy_530 <= '1';
		else
		 s_Energy_Bin_Pos_530 <= s_Energy_Bin_Pos_530;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_530 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_530;    
  
  Energy_Bin_Pos_531 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_531   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_531 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E531_C1_L_Pos and PEAK_C1_Pos <= s_E531_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_531 <= s_Energy_Bin_Pos_531 +'1';
		 Energy_Bin_Pos_Rdy_531 <= '1';
		else
		 s_Energy_Bin_Pos_531 <= s_Energy_Bin_Pos_531;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_531 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_531;   
  
  Energy_Bin_Pos_532 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_532   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_532 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E532_C1_L_Pos and PEAK_C1_Pos <= s_E532_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_532 <= s_Energy_Bin_Pos_532 +'1';
		 Energy_Bin_Pos_Rdy_532 <= '1';
		else
		 s_Energy_Bin_Pos_532 <= s_Energy_Bin_Pos_532;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_532 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_532;   
  
  Energy_Bin_Pos_533 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_533   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_533 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E533_C1_L_Pos and PEAK_C1_Pos <= s_E533_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_533 <= s_Energy_Bin_Pos_533 +'1';
		 Energy_Bin_Pos_Rdy_533 <= '1';
		else
		 s_Energy_Bin_Pos_533 <= s_Energy_Bin_Pos_533;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_533 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_533;   
  
  Energy_Bin_Pos_534 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_534   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_534 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E534_C1_L_Pos and PEAK_C1_Pos <= s_E534_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_534 <= s_Energy_Bin_Pos_534 +'1';
		 Energy_Bin_Pos_Rdy_534 <= '1';
		else
		 s_Energy_Bin_Pos_534 <= s_Energy_Bin_Pos_534;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_534 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_534;   
 
 
  Energy_Bin_Pos_535 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_535   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_535 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E535_C1_L_Pos and PEAK_C1_Pos <= s_E535_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_535 <= s_Energy_Bin_Pos_535 +'1';
		 Energy_Bin_Pos_Rdy_535 <= '1';
		else
		 s_Energy_Bin_Pos_535 <= s_Energy_Bin_Pos_535;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_535 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_535;  
 
  
  Energy_Bin_Pos_536 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_536   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_536 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E536_C1_L_Pos and PEAK_C1_Pos <= s_E536_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_536 <= s_Energy_Bin_Pos_536 +'1';
		 Energy_Bin_Pos_Rdy_536 <= '1';
		else
		 s_Energy_Bin_Pos_536 <= s_Energy_Bin_Pos_536;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_536 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_536;   
  
 Energy_Bin_Pos_537 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_537   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_537 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E537_C1_L_Pos and PEAK_C1_Pos <= s_E537_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_537 <= s_Energy_Bin_Pos_537 +'1';
		 Energy_Bin_Pos_Rdy_537 <= '1';
		else
		 s_Energy_Bin_Pos_537 <= s_Energy_Bin_Pos_537;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_537 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_537;   
  
  Energy_Bin_Pos_538 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_538   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_538 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E538_C1_L_Pos and PEAK_C1_Pos <= s_E538_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_538 <= s_Energy_Bin_Pos_538 +'1';
		 Energy_Bin_Pos_Rdy_538 <= '1';
		else
		 s_Energy_Bin_Pos_538 <= s_Energy_Bin_Pos_538;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_538 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_538;   
  
  Energy_Bin_Pos_539 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_539   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_539 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E539_C1_L_Pos and PEAK_C1_Pos <= s_E539_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_539 <= s_Energy_Bin_Pos_539 +'1';
		 Energy_Bin_Pos_Rdy_539 <= '1';
		else
		 s_Energy_Bin_Pos_539 <= s_Energy_Bin_Pos_539;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_539 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_539;         
  
     Energy_Bin_Pos_540 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_540   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_540 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E540_C1_L_Pos and PEAK_C1_Pos <= s_E540_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_540 <= s_Energy_Bin_Pos_540 +'1';
		 Energy_Bin_Pos_Rdy_540 <= '1';
		else
		 s_Energy_Bin_Pos_540 <= s_Energy_Bin_Pos_540;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_540 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_540;    
  
  Energy_Bin_Pos_541 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_541   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_541 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E541_C1_L_Pos and PEAK_C1_Pos <= s_E541_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_541 <= s_Energy_Bin_Pos_541 +'1';
		 Energy_Bin_Pos_Rdy_541 <= '1';
		else
		 s_Energy_Bin_Pos_541 <= s_Energy_Bin_Pos_541;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_541 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_541;   
  
  Energy_Bin_Pos_542 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_542   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_542 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E542_C1_L_Pos and PEAK_C1_Pos <= s_E542_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_542 <= s_Energy_Bin_Pos_542 +'1';
		 Energy_Bin_Pos_Rdy_542 <= '1';
		else
		 s_Energy_Bin_Pos_542 <= s_Energy_Bin_Pos_542;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_542 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_542;   
  
  Energy_Bin_Pos_543 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_543   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_543 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E543_C1_L_Pos and PEAK_C1_Pos <= s_E543_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_543 <= s_Energy_Bin_Pos_543 +'1';
		 Energy_Bin_Pos_Rdy_543 <= '1';
		else
		 s_Energy_Bin_Pos_543 <= s_Energy_Bin_Pos_543;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_543 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_543;   
  
  Energy_Bin_Pos_544 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_544   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_544 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E544_C1_L_Pos and PEAK_C1_Pos <= s_E544_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_544 <= s_Energy_Bin_Pos_544 +'1';
		 Energy_Bin_Pos_Rdy_544 <= '1';
		else
		 s_Energy_Bin_Pos_544 <= s_Energy_Bin_Pos_544;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_544 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_544;   
 
 
  Energy_Bin_Pos_545 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_545   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_545 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E545_C1_L_Pos and PEAK_C1_Pos <= s_E545_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_545 <= s_Energy_Bin_Pos_545 +'1';
		 Energy_Bin_Pos_Rdy_545 <= '1';
		else
		 s_Energy_Bin_Pos_545 <= s_Energy_Bin_Pos_545;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_545 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_545;  
 
  
  Energy_Bin_Pos_546 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_546   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_546 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E546_C1_L_Pos and PEAK_C1_Pos <= s_E546_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_546 <= s_Energy_Bin_Pos_546 +'1';
		 Energy_Bin_Pos_Rdy_546 <= '1';
		else
		 s_Energy_Bin_Pos_546 <= s_Energy_Bin_Pos_546;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_546 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_546;   
  
 Energy_Bin_Pos_547 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_547   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_547 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E547_C1_L_Pos and PEAK_C1_Pos <= s_E547_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_547 <= s_Energy_Bin_Pos_547 +'1';
		 Energy_Bin_Pos_Rdy_547 <= '1';
		else
		 s_Energy_Bin_Pos_547 <= s_Energy_Bin_Pos_547;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_547 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_547;   
  
  Energy_Bin_Pos_548 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_548   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_548 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E548_C1_L_Pos and PEAK_C1_Pos <= s_E548_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_548 <= s_Energy_Bin_Pos_548 +'1';
		 Energy_Bin_Pos_Rdy_548 <= '1';
		else
		 s_Energy_Bin_Pos_548 <= s_Energy_Bin_Pos_548;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_548 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_548;   
  
  Energy_Bin_Pos_549 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_549   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_549 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E549_C1_L_Pos and PEAK_C1_Pos <= s_E549_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_549 <= s_Energy_Bin_Pos_549 +'1';
		 Energy_Bin_Pos_Rdy_549 <= '1';
		else
		 s_Energy_Bin_Pos_549 <= s_Energy_Bin_Pos_549;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_549 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_549;          
  
  
     Energy_Bin_Pos_550 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_550   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_550 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E550_C1_L_Pos and PEAK_C1_Pos <= s_E550_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_550 <= s_Energy_Bin_Pos_550 +'1';
		 Energy_Bin_Pos_Rdy_550 <= '1';
		else
		 s_Energy_Bin_Pos_550 <= s_Energy_Bin_Pos_550;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_550 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_550;    
  
  Energy_Bin_Pos_551 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_551   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_551 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E551_C1_L_Pos and PEAK_C1_Pos <= s_E551_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_551 <= s_Energy_Bin_Pos_551 +'1';
		 Energy_Bin_Pos_Rdy_551 <= '1';
		else
		 s_Energy_Bin_Pos_551 <= s_Energy_Bin_Pos_551;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_551 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_551;   
  
  Energy_Bin_Pos_552 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_552   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_552 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E552_C1_L_Pos and PEAK_C1_Pos <= s_E552_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_552 <= s_Energy_Bin_Pos_552 +'1';
		 Energy_Bin_Pos_Rdy_552 <= '1';
		else
		 s_Energy_Bin_Pos_552 <= s_Energy_Bin_Pos_552;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_552 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_552;   
  
  Energy_Bin_Pos_553 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_553   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_553 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E553_C1_L_Pos and PEAK_C1_Pos <= s_E553_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_553 <= s_Energy_Bin_Pos_553 +'1';
		 Energy_Bin_Pos_Rdy_553 <= '1';
		else
		 s_Energy_Bin_Pos_553 <= s_Energy_Bin_Pos_553;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_553 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_553;   
  
  Energy_Bin_Pos_554 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_554   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_554 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E554_C1_L_Pos and PEAK_C1_Pos <= s_E554_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_554 <= s_Energy_Bin_Pos_554 +'1';
		 Energy_Bin_Pos_Rdy_554 <= '1';
		else
		 s_Energy_Bin_Pos_554 <= s_Energy_Bin_Pos_554;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_554 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_554;   
 
 
  Energy_Bin_Pos_555 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_555   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_555 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E555_C1_L_Pos and PEAK_C1_Pos <= s_E555_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_555 <= s_Energy_Bin_Pos_555 +'1';
		 Energy_Bin_Pos_Rdy_555 <= '1';
		else
		 s_Energy_Bin_Pos_555 <= s_Energy_Bin_Pos_555;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_555 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_555;  
 
  
  Energy_Bin_Pos_556 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_556   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_556 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E556_C1_L_Pos and PEAK_C1_Pos <= s_E556_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_556 <= s_Energy_Bin_Pos_556 +'1';
		 Energy_Bin_Pos_Rdy_556 <= '1';
		else
		 s_Energy_Bin_Pos_556 <= s_Energy_Bin_Pos_556;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_556 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_556;   
  
 Energy_Bin_Pos_557 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_557   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_557 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E557_C1_L_Pos and PEAK_C1_Pos <= s_E557_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_557 <= s_Energy_Bin_Pos_557 +'1';
		 Energy_Bin_Pos_Rdy_557 <= '1';
		else
		 s_Energy_Bin_Pos_557 <= s_Energy_Bin_Pos_557;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_557 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_557;   
  
  Energy_Bin_Pos_558 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_558   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_558 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E558_C1_L_Pos and PEAK_C1_Pos <= s_E558_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_558 <= s_Energy_Bin_Pos_558 +'1';
		 Energy_Bin_Pos_Rdy_558 <= '1';
		else
		 s_Energy_Bin_Pos_558 <= s_Energy_Bin_Pos_558;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_558 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_558;   
  
  Energy_Bin_Pos_559 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_559   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_559 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E559_C1_L_Pos and PEAK_C1_Pos <= s_E559_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_559 <= s_Energy_Bin_Pos_559 +'1';
		 Energy_Bin_Pos_Rdy_559 <= '1';
		else
		 s_Energy_Bin_Pos_559 <= s_Energy_Bin_Pos_559;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_559 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_559;           
  
     Energy_Bin_Pos_560 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_560   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_560 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E560_C1_L_Pos and PEAK_C1_Pos <= s_E560_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_560 <= s_Energy_Bin_Pos_560 +'1';
		 Energy_Bin_Pos_Rdy_560 <= '1';
		else
		 s_Energy_Bin_Pos_560 <= s_Energy_Bin_Pos_560;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_560 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_560;    
  
  Energy_Bin_Pos_561 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_561   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_561 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E561_C1_L_Pos and PEAK_C1_Pos <= s_E561_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_561 <= s_Energy_Bin_Pos_561 +'1';
		 Energy_Bin_Pos_Rdy_561 <= '1';
		else
		 s_Energy_Bin_Pos_561 <= s_Energy_Bin_Pos_561;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_561 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_561;   
  
  Energy_Bin_Pos_562 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_562   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_562 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E562_C1_L_Pos and PEAK_C1_Pos <= s_E562_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_562 <= s_Energy_Bin_Pos_562 +'1';
		 Energy_Bin_Pos_Rdy_562 <= '1';
		else
		 s_Energy_Bin_Pos_562 <= s_Energy_Bin_Pos_562;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_562 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_562;   
  
  Energy_Bin_Pos_563 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_563   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_563 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E563_C1_L_Pos and PEAK_C1_Pos <= s_E563_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_563 <= s_Energy_Bin_Pos_563 +'1';
		 Energy_Bin_Pos_Rdy_563 <= '1';
		else
		 s_Energy_Bin_Pos_563 <= s_Energy_Bin_Pos_563;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_563 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_563;   
  
  Energy_Bin_Pos_564 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_564   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_564 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E564_C1_L_Pos and PEAK_C1_Pos <= s_E564_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_564 <= s_Energy_Bin_Pos_564 +'1';
		 Energy_Bin_Pos_Rdy_564 <= '1';
		else
		 s_Energy_Bin_Pos_564 <= s_Energy_Bin_Pos_564;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_564 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_564;   
 
 
  Energy_Bin_Pos_565 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_565   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_565 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E565_C1_L_Pos and PEAK_C1_Pos <= s_E565_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_565 <= s_Energy_Bin_Pos_565 +'1';
		 Energy_Bin_Pos_Rdy_565 <= '1';
		else
		 s_Energy_Bin_Pos_565 <= s_Energy_Bin_Pos_565;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_565 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_565;  
 
  
  Energy_Bin_Pos_566 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_566   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_566 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E566_C1_L_Pos and PEAK_C1_Pos <= s_E566_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_566 <= s_Energy_Bin_Pos_566 +'1';
		 Energy_Bin_Pos_Rdy_566 <= '1';
		else
		 s_Energy_Bin_Pos_566 <= s_Energy_Bin_Pos_566;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_566 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_566;   
  
 Energy_Bin_Pos_567 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_567   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_567 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E567_C1_L_Pos and PEAK_C1_Pos <= s_E567_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_567 <= s_Energy_Bin_Pos_567 +'1';
		 Energy_Bin_Pos_Rdy_567 <= '1';
		else
		 s_Energy_Bin_Pos_567 <= s_Energy_Bin_Pos_567;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_567 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_567;   
  
  Energy_Bin_Pos_568 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_568   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_568 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E568_C1_L_Pos and PEAK_C1_Pos <= s_E568_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_568 <= s_Energy_Bin_Pos_568 +'1';
		 Energy_Bin_Pos_Rdy_568 <= '1';
		else
		 s_Energy_Bin_Pos_568 <= s_Energy_Bin_Pos_568;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_568 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_568;   
  
  Energy_Bin_Pos_569 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_569   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_569 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E569_C1_L_Pos and PEAK_C1_Pos <= s_E569_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_569 <= s_Energy_Bin_Pos_569 +'1';
		 Energy_Bin_Pos_Rdy_569 <= '1';
		else
		 s_Energy_Bin_Pos_569 <= s_Energy_Bin_Pos_569;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_569 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_569;         
  
     Energy_Bin_Pos_570 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_570   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_570 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E570_C1_L_Pos and PEAK_C1_Pos <= s_E570_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_570 <= s_Energy_Bin_Pos_570 +'1';
		 Energy_Bin_Pos_Rdy_570 <= '1';
		else
		 s_Energy_Bin_Pos_570 <= s_Energy_Bin_Pos_570;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_570 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_570;    
  
  Energy_Bin_Pos_571 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_571   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_571 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E571_C1_L_Pos and PEAK_C1_Pos <= s_E571_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_571 <= s_Energy_Bin_Pos_571 +'1';
		 Energy_Bin_Pos_Rdy_571 <= '1';
		else
		 s_Energy_Bin_Pos_571 <= s_Energy_Bin_Pos_571;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_571 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_571;   
  
  Energy_Bin_Pos_572 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_572   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_572 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E572_C1_L_Pos and PEAK_C1_Pos <= s_E572_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_572 <= s_Energy_Bin_Pos_572 +'1';
		 Energy_Bin_Pos_Rdy_572 <= '1';
		else
		 s_Energy_Bin_Pos_572 <= s_Energy_Bin_Pos_572;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_572 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_572;   
  
  Energy_Bin_Pos_573 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_573   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_573 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E573_C1_L_Pos and PEAK_C1_Pos <= s_E573_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_573 <= s_Energy_Bin_Pos_573 +'1';
		 Energy_Bin_Pos_Rdy_573 <= '1';
		else
		 s_Energy_Bin_Pos_573 <= s_Energy_Bin_Pos_573;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_573 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_573;   
  
  Energy_Bin_Pos_574 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_574   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_574 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E574_C1_L_Pos and PEAK_C1_Pos <= s_E574_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_574 <= s_Energy_Bin_Pos_574 +'1';
		 Energy_Bin_Pos_Rdy_574 <= '1';
		else
		 s_Energy_Bin_Pos_574 <= s_Energy_Bin_Pos_574;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_574 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_574;   
 
 
  Energy_Bin_Pos_575 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_575   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_575 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E575_C1_L_Pos and PEAK_C1_Pos <= s_E575_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_575 <= s_Energy_Bin_Pos_575 +'1';
		 Energy_Bin_Pos_Rdy_575 <= '1';
		else
		 s_Energy_Bin_Pos_575 <= s_Energy_Bin_Pos_575;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_575 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_575;  
 
  
  Energy_Bin_Pos_576 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_576   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_576 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E576_C1_L_Pos and PEAK_C1_Pos <= s_E576_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_576 <= s_Energy_Bin_Pos_576 +'1';
		 Energy_Bin_Pos_Rdy_576 <= '1';
		else
		 s_Energy_Bin_Pos_576 <= s_Energy_Bin_Pos_576;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_576 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_576;   
  
 Energy_Bin_Pos_577 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_577   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_577 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E577_C1_L_Pos and PEAK_C1_Pos <= s_E577_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_577 <= s_Energy_Bin_Pos_577 +'1';
		 Energy_Bin_Pos_Rdy_577 <= '1';
		else
		 s_Energy_Bin_Pos_577 <= s_Energy_Bin_Pos_577;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_577 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_577;   
  
  Energy_Bin_Pos_578 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_578   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_578 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E578_C1_L_Pos and PEAK_C1_Pos <= s_E578_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_578 <= s_Energy_Bin_Pos_578 +'1';
		 Energy_Bin_Pos_Rdy_578 <= '1';
		else
		 s_Energy_Bin_Pos_578 <= s_Energy_Bin_Pos_578;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_578 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_578;   
  
  Energy_Bin_Pos_579 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_579   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_579 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E579_C1_L_Pos and PEAK_C1_Pos <= s_E579_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_579 <= s_Energy_Bin_Pos_579 +'1';
		 Energy_Bin_Pos_Rdy_579 <= '1';
		else
		 s_Energy_Bin_Pos_579 <= s_Energy_Bin_Pos_579;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_579 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_579;       
  
     Energy_Bin_Pos_580 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_580   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_580 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E580_C1_L_Pos and PEAK_C1_Pos <= s_E580_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_580 <= s_Energy_Bin_Pos_580 +'1';
		 Energy_Bin_Pos_Rdy_580 <= '1';
		else
		 s_Energy_Bin_Pos_580 <= s_Energy_Bin_Pos_580;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_580 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_580;    
  
  Energy_Bin_Pos_581 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_581   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_581 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E581_C1_L_Pos and PEAK_C1_Pos <= s_E581_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_581 <= s_Energy_Bin_Pos_581 +'1';
		 Energy_Bin_Pos_Rdy_581 <= '1';
		else
		 s_Energy_Bin_Pos_581 <= s_Energy_Bin_Pos_581;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_581 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_581;   
  
  Energy_Bin_Pos_582 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_582   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_582 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E582_C1_L_Pos and PEAK_C1_Pos <= s_E582_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_582 <= s_Energy_Bin_Pos_582 +'1';
		 Energy_Bin_Pos_Rdy_582 <= '1';
		else
		 s_Energy_Bin_Pos_582 <= s_Energy_Bin_Pos_582;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_582 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_582;   
  
  Energy_Bin_Pos_583 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_583   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_583 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E583_C1_L_Pos and PEAK_C1_Pos <= s_E583_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_583 <= s_Energy_Bin_Pos_583 +'1';
		 Energy_Bin_Pos_Rdy_583 <= '1';
		else
		 s_Energy_Bin_Pos_583 <= s_Energy_Bin_Pos_583;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_583 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_583;   
  
  Energy_Bin_Pos_584 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_584   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_584 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E584_C1_L_Pos and PEAK_C1_Pos <= s_E584_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_584 <= s_Energy_Bin_Pos_584 +'1';
		 Energy_Bin_Pos_Rdy_584 <= '1';
		else
		 s_Energy_Bin_Pos_584 <= s_Energy_Bin_Pos_584;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_584 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_584;   
 
 
  Energy_Bin_Pos_585 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_585   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_585 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E585_C1_L_Pos and PEAK_C1_Pos <= s_E585_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_585 <= s_Energy_Bin_Pos_585 +'1';
		 Energy_Bin_Pos_Rdy_585 <= '1';
		else
		 s_Energy_Bin_Pos_585 <= s_Energy_Bin_Pos_585;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_585 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_585;  
 
  
  Energy_Bin_Pos_586 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_586   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_586 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E586_C1_L_Pos and PEAK_C1_Pos <= s_E586_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_586 <= s_Energy_Bin_Pos_586 +'1';
		 Energy_Bin_Pos_Rdy_586 <= '1';
		else
		 s_Energy_Bin_Pos_586 <= s_Energy_Bin_Pos_586;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_586 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_586;   
  
 Energy_Bin_Pos_587 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_587   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_587 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E587_C1_L_Pos and PEAK_C1_Pos <= s_E587_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_587 <= s_Energy_Bin_Pos_587 +'1';
		 Energy_Bin_Pos_Rdy_587 <= '1';
		else
		 s_Energy_Bin_Pos_587 <= s_Energy_Bin_Pos_587;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_587 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_587;   
  
  Energy_Bin_Pos_588 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_588   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_588 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E588_C1_L_Pos and PEAK_C1_Pos <= s_E588_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_588 <= s_Energy_Bin_Pos_588 +'1';
		 Energy_Bin_Pos_Rdy_588 <= '1';
		else
		 s_Energy_Bin_Pos_588 <= s_Energy_Bin_Pos_588;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_588 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_588;   
  
  Energy_Bin_Pos_589 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_589   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_589 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E589_C1_L_Pos and PEAK_C1_Pos <= s_E589_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_589 <= s_Energy_Bin_Pos_589 +'1';
		 Energy_Bin_Pos_Rdy_589 <= '1';
		else
		 s_Energy_Bin_Pos_589 <= s_Energy_Bin_Pos_589;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_589 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_589;      
  
     Energy_Bin_Pos_590 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_590   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_590 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E590_C1_L_Pos and PEAK_C1_Pos <= s_E590_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_590 <= s_Energy_Bin_Pos_590 +'1';
		 Energy_Bin_Pos_Rdy_590 <= '1';
		else
		 s_Energy_Bin_Pos_590 <= s_Energy_Bin_Pos_590;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_590 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_590;    
  
  Energy_Bin_Pos_591 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_591   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_591 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E591_C1_L_Pos and PEAK_C1_Pos <= s_E591_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_591 <= s_Energy_Bin_Pos_591 +'1';
		 Energy_Bin_Pos_Rdy_591 <= '1';
		else
		 s_Energy_Bin_Pos_591 <= s_Energy_Bin_Pos_591;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_591 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_591;   
  
  Energy_Bin_Pos_592 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_592   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_592 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E592_C1_L_Pos and PEAK_C1_Pos <= s_E592_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_592 <= s_Energy_Bin_Pos_592 +'1';
		 Energy_Bin_Pos_Rdy_592 <= '1';
		else
		 s_Energy_Bin_Pos_592 <= s_Energy_Bin_Pos_592;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_592 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_592;   
  
  Energy_Bin_Pos_593 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_593   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_593 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E593_C1_L_Pos and PEAK_C1_Pos <= s_E593_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_593 <= s_Energy_Bin_Pos_593 +'1';
		 Energy_Bin_Pos_Rdy_593 <= '1';
		else
		 s_Energy_Bin_Pos_593 <= s_Energy_Bin_Pos_593;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_593 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_593;   
  
  Energy_Bin_Pos_594 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_594   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_594 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E594_C1_L_Pos and PEAK_C1_Pos <= s_E594_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_594 <= s_Energy_Bin_Pos_594 +'1';
		 Energy_Bin_Pos_Rdy_594 <= '1';
		else
		 s_Energy_Bin_Pos_594 <= s_Energy_Bin_Pos_594;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_594 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_594;   
 
 
  Energy_Bin_Pos_595 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_595   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_595 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E595_C1_L_Pos and PEAK_C1_Pos <= s_E595_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_595 <= s_Energy_Bin_Pos_595 +'1';
		 Energy_Bin_Pos_Rdy_595 <= '1';
		else
		 s_Energy_Bin_Pos_595 <= s_Energy_Bin_Pos_595;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_595 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_595;  
 
  
  Energy_Bin_Pos_596 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_596   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_596 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E596_C1_L_Pos and PEAK_C1_Pos <= s_E596_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_596 <= s_Energy_Bin_Pos_596 +'1';
		 Energy_Bin_Pos_Rdy_596 <= '1';
		else
		 s_Energy_Bin_Pos_596 <= s_Energy_Bin_Pos_596;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_596 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_596;   
  
 Energy_Bin_Pos_597 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_597   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_597 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E597_C1_L_Pos and PEAK_C1_Pos <= s_E597_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_597 <= s_Energy_Bin_Pos_597 +'1';
		 Energy_Bin_Pos_Rdy_597 <= '1';
		else
		 s_Energy_Bin_Pos_597 <= s_Energy_Bin_Pos_597;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_597 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_597;   
  
  Energy_Bin_Pos_598 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_598   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_598 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E598_C1_L_Pos and PEAK_C1_Pos <= s_E598_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_598 <= s_Energy_Bin_Pos_598 +'1';
		 Energy_Bin_Pos_Rdy_598 <= '1';
		else
		 s_Energy_Bin_Pos_598 <= s_Energy_Bin_Pos_598;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_598 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_598;   
  
  Energy_Bin_Pos_599 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_599   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_599 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E599_C1_L_Pos and PEAK_C1_Pos <= s_E599_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_599 <= s_Energy_Bin_Pos_599 +'1';
		 Energy_Bin_Pos_Rdy_599 <= '1';
		else
		 s_Energy_Bin_Pos_599 <= s_Energy_Bin_Pos_599;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_599 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_599;      

    Energy_Bin_Pos_600 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_600   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_600 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E600_C1_L_Pos and PEAK_C1_Pos <= s_E600_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_600 <= s_Energy_Bin_Pos_600 +'1';
		 Energy_Bin_Pos_Rdy_600 <= '1';
		else
		 s_Energy_Bin_Pos_600 <= s_Energy_Bin_Pos_600;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_600 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_600;    
  
  Energy_Bin_Pos_601 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_601   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_601 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E601_C1_L_Pos and PEAK_C1_Pos <= s_E601_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_601 <= s_Energy_Bin_Pos_601 +'1';
		 Energy_Bin_Pos_Rdy_601 <= '1';
		else
		 s_Energy_Bin_Pos_601 <= s_Energy_Bin_Pos_601;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_601 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_601;   
  
  Energy_Bin_Pos_602 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_602   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_602 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E602_C1_L_Pos and PEAK_C1_Pos <= s_E602_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_602 <= s_Energy_Bin_Pos_602 +'1';
		 Energy_Bin_Pos_Rdy_602 <= '1';
		else
		 s_Energy_Bin_Pos_602 <= s_Energy_Bin_Pos_602;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_602 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_602;   
  
  Energy_Bin_Pos_603 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_603   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_603 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E603_C1_L_Pos and PEAK_C1_Pos <= s_E603_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_603 <= s_Energy_Bin_Pos_603 +'1';
		 Energy_Bin_Pos_Rdy_603 <= '1';
		else
		 s_Energy_Bin_Pos_603 <= s_Energy_Bin_Pos_603;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_603 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_603;   
  
  Energy_Bin_Pos_604 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_604   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_604 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E604_C1_L_Pos and PEAK_C1_Pos <= s_E604_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_604 <= s_Energy_Bin_Pos_604 +'1';
		 Energy_Bin_Pos_Rdy_604 <= '1';
		else
		 s_Energy_Bin_Pos_604 <= s_Energy_Bin_Pos_604;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_604 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_604;   
 
 
  Energy_Bin_Pos_605 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_605   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_605 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E605_C1_L_Pos and PEAK_C1_Pos <= s_E605_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_605 <= s_Energy_Bin_Pos_605 +'1';
		 Energy_Bin_Pos_Rdy_605 <= '1';
		else
		 s_Energy_Bin_Pos_605 <= s_Energy_Bin_Pos_605;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_605 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_605;  
 
  
  Energy_Bin_Pos_606 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_606   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_606 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E606_C1_L_Pos and PEAK_C1_Pos <= s_E606_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_606 <= s_Energy_Bin_Pos_606 +'1';
		 Energy_Bin_Pos_Rdy_606 <= '1';
		else
		 s_Energy_Bin_Pos_606 <= s_Energy_Bin_Pos_606;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_606 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_606;   
  
 Energy_Bin_Pos_607 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_607   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_607 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E607_C1_L_Pos and PEAK_C1_Pos <= s_E607_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_607 <= s_Energy_Bin_Pos_607 +'1';
		 Energy_Bin_Pos_Rdy_607 <= '1';
		else
		 s_Energy_Bin_Pos_607 <= s_Energy_Bin_Pos_607;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_607 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_607;   
  
  Energy_Bin_Pos_608 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_608   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_608 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E608_C1_L_Pos and PEAK_C1_Pos <= s_E608_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_608 <= s_Energy_Bin_Pos_608 +'1';
		 Energy_Bin_Pos_Rdy_608 <= '1';
		else
		 s_Energy_Bin_Pos_608 <= s_Energy_Bin_Pos_608;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_608 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_608;   
  
  Energy_Bin_Pos_609 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_609   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_609 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E609_C1_L_Pos and PEAK_C1_Pos <= s_E609_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_609 <= s_Energy_Bin_Pos_609 +'1';
		 Energy_Bin_Pos_Rdy_609 <= '1';
		else
		 s_Energy_Bin_Pos_609 <= s_Energy_Bin_Pos_609;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_609 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_609;      
  
     Energy_Bin_Pos_610 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_610   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_610 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E610_C1_L_Pos and PEAK_C1_Pos <= s_E610_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_610 <= s_Energy_Bin_Pos_610 +'1';
		 Energy_Bin_Pos_Rdy_610 <= '1';
		else
		 s_Energy_Bin_Pos_610 <= s_Energy_Bin_Pos_610;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_610 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_610;    
  
  Energy_Bin_Pos_611 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_611   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_611 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E611_C1_L_Pos and PEAK_C1_Pos <= s_E611_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_611 <= s_Energy_Bin_Pos_611 +'1';
		 Energy_Bin_Pos_Rdy_611 <= '1';
		else
		 s_Energy_Bin_Pos_611 <= s_Energy_Bin_Pos_611;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_611 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_611;   
  
  Energy_Bin_Pos_612 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_612   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_612 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E612_C1_L_Pos and PEAK_C1_Pos <= s_E612_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_612 <= s_Energy_Bin_Pos_612 +'1';
		 Energy_Bin_Pos_Rdy_612 <= '1';
		else
		 s_Energy_Bin_Pos_612 <= s_Energy_Bin_Pos_612;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_612 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_612;   
  
  Energy_Bin_Pos_613 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_613   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_613 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E613_C1_L_Pos and PEAK_C1_Pos <= s_E613_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_613 <= s_Energy_Bin_Pos_613 +'1';
		 Energy_Bin_Pos_Rdy_613 <= '1';
		else
		 s_Energy_Bin_Pos_613 <= s_Energy_Bin_Pos_613;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_613 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_613;   
  
  Energy_Bin_Pos_614 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_614   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_614 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E614_C1_L_Pos and PEAK_C1_Pos <= s_E614_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_614 <= s_Energy_Bin_Pos_614 +'1';
		 Energy_Bin_Pos_Rdy_614 <= '1';
		else
		 s_Energy_Bin_Pos_614 <= s_Energy_Bin_Pos_614;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_614 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_614;   
 
 
  Energy_Bin_Pos_615 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_615   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_615 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E615_C1_L_Pos and PEAK_C1_Pos <= s_E615_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_615 <= s_Energy_Bin_Pos_615 +'1';
		 Energy_Bin_Pos_Rdy_615 <= '1';
		else
		 s_Energy_Bin_Pos_615 <= s_Energy_Bin_Pos_615;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_615 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_615;  
 
  
  Energy_Bin_Pos_616 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_616   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_616 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E616_C1_L_Pos and PEAK_C1_Pos <= s_E616_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_616 <= s_Energy_Bin_Pos_616 +'1';
		 Energy_Bin_Pos_Rdy_616 <= '1';
		else
		 s_Energy_Bin_Pos_616 <= s_Energy_Bin_Pos_616;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_616 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_616;   
  
 Energy_Bin_Pos_617 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_617   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_617 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E617_C1_L_Pos and PEAK_C1_Pos <= s_E617_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_617 <= s_Energy_Bin_Pos_617 +'1';
		 Energy_Bin_Pos_Rdy_617 <= '1';
		else
		 s_Energy_Bin_Pos_617 <= s_Energy_Bin_Pos_617;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_617 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_617;   
  
  Energy_Bin_Pos_618 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_618   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_618 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E618_C1_L_Pos and PEAK_C1_Pos <= s_E618_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_618 <= s_Energy_Bin_Pos_618 +'1';
		 Energy_Bin_Pos_Rdy_618 <= '1';
		else
		 s_Energy_Bin_Pos_618 <= s_Energy_Bin_Pos_618;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_618 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_618;   
  
  Energy_Bin_Pos_619 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_619   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_619 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E619_C1_L_Pos and PEAK_C1_Pos <= s_E619_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_619 <= s_Energy_Bin_Pos_619 +'1';
		 Energy_Bin_Pos_Rdy_619 <= '1';
		else
		 s_Energy_Bin_Pos_619 <= s_Energy_Bin_Pos_619;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_619 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_619;       
  
     Energy_Bin_Pos_620 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_620   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_620 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E620_C1_L_Pos and PEAK_C1_Pos <= s_E620_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_620 <= s_Energy_Bin_Pos_620 +'1';
		 Energy_Bin_Pos_Rdy_620 <= '1';
		else
		 s_Energy_Bin_Pos_620 <= s_Energy_Bin_Pos_620;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_620 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_620;    
  
  Energy_Bin_Pos_621 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_621   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_621 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E621_C1_L_Pos and PEAK_C1_Pos <= s_E621_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_621 <= s_Energy_Bin_Pos_621 +'1';
		 Energy_Bin_Pos_Rdy_621 <= '1';
		else
		 s_Energy_Bin_Pos_621 <= s_Energy_Bin_Pos_621;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_621 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_621;   
  
  Energy_Bin_Pos_622 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_622   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_622 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E622_C1_L_Pos and PEAK_C1_Pos <= s_E622_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_622 <= s_Energy_Bin_Pos_622 +'1';
		 Energy_Bin_Pos_Rdy_622 <= '1';
		else
		 s_Energy_Bin_Pos_622 <= s_Energy_Bin_Pos_622;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_622 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_622;   
  
  Energy_Bin_Pos_623 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_623   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_623 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E623_C1_L_Pos and PEAK_C1_Pos <= s_E623_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_623 <= s_Energy_Bin_Pos_623 +'1';
		 Energy_Bin_Pos_Rdy_623 <= '1';
		else
		 s_Energy_Bin_Pos_623 <= s_Energy_Bin_Pos_623;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_623 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_623;   
  
  Energy_Bin_Pos_624 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_624   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_624 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E624_C1_L_Pos and PEAK_C1_Pos <= s_E624_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_624 <= s_Energy_Bin_Pos_624 +'1';
		 Energy_Bin_Pos_Rdy_624 <= '1';
		else
		 s_Energy_Bin_Pos_624 <= s_Energy_Bin_Pos_624;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_624 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_624;   
 
 
  Energy_Bin_Pos_625 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_625   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_625 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E625_C1_L_Pos and PEAK_C1_Pos <= s_E625_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_625 <= s_Energy_Bin_Pos_625 +'1';
		 Energy_Bin_Pos_Rdy_625 <= '1';
		else
		 s_Energy_Bin_Pos_625 <= s_Energy_Bin_Pos_625;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_625 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_625;  
 
  
  Energy_Bin_Pos_626 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_626   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_626 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E626_C1_L_Pos and PEAK_C1_Pos <= s_E626_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_626 <= s_Energy_Bin_Pos_626 +'1';
		 Energy_Bin_Pos_Rdy_626 <= '1';
		else
		 s_Energy_Bin_Pos_626 <= s_Energy_Bin_Pos_626;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_626 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_626;   
  
 Energy_Bin_Pos_627 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_627   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_627 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E627_C1_L_Pos and PEAK_C1_Pos <= s_E627_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_627 <= s_Energy_Bin_Pos_627 +'1';
		 Energy_Bin_Pos_Rdy_627 <= '1';
		else
		 s_Energy_Bin_Pos_627 <= s_Energy_Bin_Pos_627;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_627 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_627;   
  
  Energy_Bin_Pos_628 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_628   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_628 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E628_C1_L_Pos and PEAK_C1_Pos <= s_E628_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_628 <= s_Energy_Bin_Pos_628 +'1';
		 Energy_Bin_Pos_Rdy_628 <= '1';
		else
		 s_Energy_Bin_Pos_628 <= s_Energy_Bin_Pos_628;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_628 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_628;   
  
  Energy_Bin_Pos_629 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_629   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_629 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E629_C1_L_Pos and PEAK_C1_Pos <= s_E629_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_629 <= s_Energy_Bin_Pos_629 +'1';
		 Energy_Bin_Pos_Rdy_629 <= '1';
		else
		 s_Energy_Bin_Pos_629 <= s_Energy_Bin_Pos_629;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_629 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_629;        
  
     Energy_Bin_Pos_630 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_630   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_630 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E630_C1_L_Pos and PEAK_C1_Pos <= s_E630_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_630 <= s_Energy_Bin_Pos_630 +'1';
		 Energy_Bin_Pos_Rdy_630 <= '1';
		else
		 s_Energy_Bin_Pos_630 <= s_Energy_Bin_Pos_630;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_630 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_630;    
  
  Energy_Bin_Pos_631 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_631   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_631 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E631_C1_L_Pos and PEAK_C1_Pos <= s_E631_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_631 <= s_Energy_Bin_Pos_631 +'1';
		 Energy_Bin_Pos_Rdy_631 <= '1';
		else
		 s_Energy_Bin_Pos_631 <= s_Energy_Bin_Pos_631;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_631 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_631;   
  
  Energy_Bin_Pos_632 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_632   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_632 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E632_C1_L_Pos and PEAK_C1_Pos <= s_E632_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_632 <= s_Energy_Bin_Pos_632 +'1';
		 Energy_Bin_Pos_Rdy_632 <= '1';
		else
		 s_Energy_Bin_Pos_632 <= s_Energy_Bin_Pos_632;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_632 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_632;   
  
  Energy_Bin_Pos_633 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_633   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_633 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E633_C1_L_Pos and PEAK_C1_Pos <= s_E633_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_633 <= s_Energy_Bin_Pos_633 +'1';
		 Energy_Bin_Pos_Rdy_633 <= '1';
		else
		 s_Energy_Bin_Pos_633 <= s_Energy_Bin_Pos_633;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_633 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_633;   
  
  Energy_Bin_Pos_634 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_634   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_634 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E634_C1_L_Pos and PEAK_C1_Pos <= s_E634_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_634 <= s_Energy_Bin_Pos_634 +'1';
		 Energy_Bin_Pos_Rdy_634 <= '1';
		else
		 s_Energy_Bin_Pos_634 <= s_Energy_Bin_Pos_634;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_634 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_634;   
 
 
  Energy_Bin_Pos_635 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_635   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_635 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E635_C1_L_Pos and PEAK_C1_Pos <= s_E635_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_635 <= s_Energy_Bin_Pos_635 +'1';
		 Energy_Bin_Pos_Rdy_635 <= '1';
		else
		 s_Energy_Bin_Pos_635 <= s_Energy_Bin_Pos_635;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_635 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_635;  
 
  
  Energy_Bin_Pos_636 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_636   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_636 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E636_C1_L_Pos and PEAK_C1_Pos <= s_E636_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_636 <= s_Energy_Bin_Pos_636 +'1';
		 Energy_Bin_Pos_Rdy_636 <= '1';
		else
		 s_Energy_Bin_Pos_636 <= s_Energy_Bin_Pos_636;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_636 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_636;   
  
 Energy_Bin_Pos_637 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_637   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_637 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E637_C1_L_Pos and PEAK_C1_Pos <= s_E637_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_637 <= s_Energy_Bin_Pos_637 +'1';
		 Energy_Bin_Pos_Rdy_637 <= '1';
		else
		 s_Energy_Bin_Pos_637 <= s_Energy_Bin_Pos_637;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_637 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_637;   
  
  Energy_Bin_Pos_638 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_638   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_638 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E638_C1_L_Pos and PEAK_C1_Pos <= s_E638_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_638 <= s_Energy_Bin_Pos_638 +'1';
		 Energy_Bin_Pos_Rdy_638 <= '1';
		else
		 s_Energy_Bin_Pos_638 <= s_Energy_Bin_Pos_638;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_638 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_638;   
  
  Energy_Bin_Pos_639 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_639   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_639 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E639_C1_L_Pos and PEAK_C1_Pos <= s_E639_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_639 <= s_Energy_Bin_Pos_639 +'1';
		 Energy_Bin_Pos_Rdy_639 <= '1';
		else
		 s_Energy_Bin_Pos_639 <= s_Energy_Bin_Pos_639;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_639 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_639;         
  
     Energy_Bin_Pos_640 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_640   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_640 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E640_C1_L_Pos and PEAK_C1_Pos <= s_E640_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_640 <= s_Energy_Bin_Pos_640 +'1';
		 Energy_Bin_Pos_Rdy_640 <= '1';
		else
		 s_Energy_Bin_Pos_640 <= s_Energy_Bin_Pos_640;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_640 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_640;    
  
  Energy_Bin_Pos_641 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_641   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_641 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E641_C1_L_Pos and PEAK_C1_Pos <= s_E641_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_641 <= s_Energy_Bin_Pos_641 +'1';
		 Energy_Bin_Pos_Rdy_641 <= '1';
		else
		 s_Energy_Bin_Pos_641 <= s_Energy_Bin_Pos_641;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_641 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_641;   
  
  Energy_Bin_Pos_642 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_642   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_642 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E642_C1_L_Pos and PEAK_C1_Pos <= s_E642_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_642 <= s_Energy_Bin_Pos_642 +'1';
		 Energy_Bin_Pos_Rdy_642 <= '1';
		else
		 s_Energy_Bin_Pos_642 <= s_Energy_Bin_Pos_642;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_642 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_642;   
  
  Energy_Bin_Pos_643 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_643   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_643 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E643_C1_L_Pos and PEAK_C1_Pos <= s_E643_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_643 <= s_Energy_Bin_Pos_643 +'1';
		 Energy_Bin_Pos_Rdy_643 <= '1';
		else
		 s_Energy_Bin_Pos_643 <= s_Energy_Bin_Pos_643;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_643 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_643;   
  
  Energy_Bin_Pos_644 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_644   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_644 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E644_C1_L_Pos and PEAK_C1_Pos <= s_E644_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_644 <= s_Energy_Bin_Pos_644 +'1';
		 Energy_Bin_Pos_Rdy_644 <= '1';
		else
		 s_Energy_Bin_Pos_644 <= s_Energy_Bin_Pos_644;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_644 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_644;   
 
 
  Energy_Bin_Pos_645 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_645   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_645 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E645_C1_L_Pos and PEAK_C1_Pos <= s_E645_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_645 <= s_Energy_Bin_Pos_645 +'1';
		 Energy_Bin_Pos_Rdy_645 <= '1';
		else
		 s_Energy_Bin_Pos_645 <= s_Energy_Bin_Pos_645;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_645 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_645;  
 
  
  Energy_Bin_Pos_646 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_646   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_646 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E646_C1_L_Pos and PEAK_C1_Pos <= s_E646_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_646 <= s_Energy_Bin_Pos_646 +'1';
		 Energy_Bin_Pos_Rdy_646 <= '1';
		else
		 s_Energy_Bin_Pos_646 <= s_Energy_Bin_Pos_646;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_646 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_646;   
  
 Energy_Bin_Pos_647 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_647   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_647 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E647_C1_L_Pos and PEAK_C1_Pos <= s_E647_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_647 <= s_Energy_Bin_Pos_647 +'1';
		 Energy_Bin_Pos_Rdy_647 <= '1';
		else
		 s_Energy_Bin_Pos_647 <= s_Energy_Bin_Pos_647;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_647 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_647;   
  
  Energy_Bin_Pos_648 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_648   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_648 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E648_C1_L_Pos and PEAK_C1_Pos <= s_E648_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_648 <= s_Energy_Bin_Pos_648 +'1';
		 Energy_Bin_Pos_Rdy_648 <= '1';
		else
		 s_Energy_Bin_Pos_648 <= s_Energy_Bin_Pos_648;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_648 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_648;   
  
  Energy_Bin_Pos_649 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_649   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_649 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E649_C1_L_Pos and PEAK_C1_Pos <= s_E649_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_649 <= s_Energy_Bin_Pos_649 +'1';
		 Energy_Bin_Pos_Rdy_649 <= '1';
		else
		 s_Energy_Bin_Pos_649 <= s_Energy_Bin_Pos_649;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_649 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_649;          
  
  
     Energy_Bin_Pos_650 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_650   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_650 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E650_C1_L_Pos and PEAK_C1_Pos <= s_E650_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_650 <= s_Energy_Bin_Pos_650 +'1';
		 Energy_Bin_Pos_Rdy_650 <= '1';
		else
		 s_Energy_Bin_Pos_650 <= s_Energy_Bin_Pos_650;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_650 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_650;    
  
  Energy_Bin_Pos_651 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_651   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_651 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E651_C1_L_Pos and PEAK_C1_Pos <= s_E651_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_651 <= s_Energy_Bin_Pos_651 +'1';
		 Energy_Bin_Pos_Rdy_651 <= '1';
		else
		 s_Energy_Bin_Pos_651 <= s_Energy_Bin_Pos_651;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_651 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_651;   
  
  Energy_Bin_Pos_652 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_652   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_652 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E652_C1_L_Pos and PEAK_C1_Pos <= s_E652_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_652 <= s_Energy_Bin_Pos_652 +'1';
		 Energy_Bin_Pos_Rdy_652 <= '1';
		else
		 s_Energy_Bin_Pos_652 <= s_Energy_Bin_Pos_652;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_652 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_652;   
  
  Energy_Bin_Pos_653 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_653   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_653 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E653_C1_L_Pos and PEAK_C1_Pos <= s_E653_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_653 <= s_Energy_Bin_Pos_653 +'1';
		 Energy_Bin_Pos_Rdy_653 <= '1';
		else
		 s_Energy_Bin_Pos_653 <= s_Energy_Bin_Pos_653;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_653 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_653;   
  
  Energy_Bin_Pos_654 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_654   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_654 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E654_C1_L_Pos and PEAK_C1_Pos <= s_E654_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_654 <= s_Energy_Bin_Pos_654 +'1';
		 Energy_Bin_Pos_Rdy_654 <= '1';
		else
		 s_Energy_Bin_Pos_654 <= s_Energy_Bin_Pos_654;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_654 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_654;   
 
 
  Energy_Bin_Pos_655 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_655   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_655 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E655_C1_L_Pos and PEAK_C1_Pos <= s_E655_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_655 <= s_Energy_Bin_Pos_655 +'1';
		 Energy_Bin_Pos_Rdy_655 <= '1';
		else
		 s_Energy_Bin_Pos_655 <= s_Energy_Bin_Pos_655;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_655 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_655;  
 
  
  Energy_Bin_Pos_656 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_656   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_656 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E656_C1_L_Pos and PEAK_C1_Pos <= s_E656_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_656 <= s_Energy_Bin_Pos_656 +'1';
		 Energy_Bin_Pos_Rdy_656 <= '1';
		else
		 s_Energy_Bin_Pos_656 <= s_Energy_Bin_Pos_656;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_656 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_656;   
  
 Energy_Bin_Pos_657 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_657   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_657 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E657_C1_L_Pos and PEAK_C1_Pos <= s_E657_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_657 <= s_Energy_Bin_Pos_657 +'1';
		 Energy_Bin_Pos_Rdy_657 <= '1';
		else
		 s_Energy_Bin_Pos_657 <= s_Energy_Bin_Pos_657;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_657 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_657;   
  
  Energy_Bin_Pos_658 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_658   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_658 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E658_C1_L_Pos and PEAK_C1_Pos <= s_E658_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_658 <= s_Energy_Bin_Pos_658 +'1';
		 Energy_Bin_Pos_Rdy_658 <= '1';
		else
		 s_Energy_Bin_Pos_658 <= s_Energy_Bin_Pos_658;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_658 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_658;   
  
  Energy_Bin_Pos_659 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_659   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_659 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E659_C1_L_Pos and PEAK_C1_Pos <= s_E659_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_659 <= s_Energy_Bin_Pos_659 +'1';
		 Energy_Bin_Pos_Rdy_659 <= '1';
		else
		 s_Energy_Bin_Pos_659 <= s_Energy_Bin_Pos_659;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_659 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_659;           
  
     Energy_Bin_Pos_660 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_660   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_660 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E660_C1_L_Pos and PEAK_C1_Pos <= s_E660_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_660 <= s_Energy_Bin_Pos_660 +'1';
		 Energy_Bin_Pos_Rdy_660 <= '1';
		else
		 s_Energy_Bin_Pos_660 <= s_Energy_Bin_Pos_660;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_660 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_660;    
  
  Energy_Bin_Pos_661 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_661   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_661 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E661_C1_L_Pos and PEAK_C1_Pos <= s_E661_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_661 <= s_Energy_Bin_Pos_661 +'1';
		 Energy_Bin_Pos_Rdy_661 <= '1';
		else
		 s_Energy_Bin_Pos_661 <= s_Energy_Bin_Pos_661;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_661 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_661;   
  
  Energy_Bin_Pos_662 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_662   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_662 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E662_C1_L_Pos and PEAK_C1_Pos <= s_E662_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_662 <= s_Energy_Bin_Pos_662 +'1';
		 Energy_Bin_Pos_Rdy_662 <= '1';
		else
		 s_Energy_Bin_Pos_662 <= s_Energy_Bin_Pos_662;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_662 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_662;   
  
  Energy_Bin_Pos_663 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_663   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_663 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E663_C1_L_Pos and PEAK_C1_Pos <= s_E663_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_663 <= s_Energy_Bin_Pos_663 +'1';
		 Energy_Bin_Pos_Rdy_663 <= '1';
		else
		 s_Energy_Bin_Pos_663 <= s_Energy_Bin_Pos_663;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_663 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_663;   
  
  Energy_Bin_Pos_664 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_664   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_664 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E664_C1_L_Pos and PEAK_C1_Pos <= s_E664_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_664 <= s_Energy_Bin_Pos_664 +'1';
		 Energy_Bin_Pos_Rdy_664 <= '1';
		else
		 s_Energy_Bin_Pos_664 <= s_Energy_Bin_Pos_664;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_664 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_664;   
 
 
  Energy_Bin_Pos_665 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_665   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_665 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E665_C1_L_Pos and PEAK_C1_Pos <= s_E665_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_665 <= s_Energy_Bin_Pos_665 +'1';
		 Energy_Bin_Pos_Rdy_665 <= '1';
		else
		 s_Energy_Bin_Pos_665 <= s_Energy_Bin_Pos_665;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_665 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_665;  
 
  
  Energy_Bin_Pos_666 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_666   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_666 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E666_C1_L_Pos and PEAK_C1_Pos <= s_E666_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_666 <= s_Energy_Bin_Pos_666 +'1';
		 Energy_Bin_Pos_Rdy_666 <= '1';
		else
		 s_Energy_Bin_Pos_666 <= s_Energy_Bin_Pos_666;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_666 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_666;   
  
 Energy_Bin_Pos_667 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_667   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_667 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E667_C1_L_Pos and PEAK_C1_Pos <= s_E667_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_667 <= s_Energy_Bin_Pos_667 +'1';
		 Energy_Bin_Pos_Rdy_667 <= '1';
		else
		 s_Energy_Bin_Pos_667 <= s_Energy_Bin_Pos_667;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_667 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_667;   
  
  Energy_Bin_Pos_668 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_668   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_668 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E668_C1_L_Pos and PEAK_C1_Pos <= s_E668_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_668 <= s_Energy_Bin_Pos_668 +'1';
		 Energy_Bin_Pos_Rdy_668 <= '1';
		else
		 s_Energy_Bin_Pos_668 <= s_Energy_Bin_Pos_668;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_668 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_668;   
  
  Energy_Bin_Pos_669 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_669   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_669 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E669_C1_L_Pos and PEAK_C1_Pos <= s_E669_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_669 <= s_Energy_Bin_Pos_669 +'1';
		 Energy_Bin_Pos_Rdy_669 <= '1';
		else
		 s_Energy_Bin_Pos_669 <= s_Energy_Bin_Pos_669;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_669 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_669;         
  
     Energy_Bin_Pos_670 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_670   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_670 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E670_C1_L_Pos and PEAK_C1_Pos <= s_E670_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_670 <= s_Energy_Bin_Pos_670 +'1';
		 Energy_Bin_Pos_Rdy_670 <= '1';
		else
		 s_Energy_Bin_Pos_670 <= s_Energy_Bin_Pos_670;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_670 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_670;    
  
  Energy_Bin_Pos_671 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_671   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_671 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E671_C1_L_Pos and PEAK_C1_Pos <= s_E671_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_671 <= s_Energy_Bin_Pos_671 +'1';
		 Energy_Bin_Pos_Rdy_671 <= '1';
		else
		 s_Energy_Bin_Pos_671 <= s_Energy_Bin_Pos_671;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_671 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_671;   
  
  Energy_Bin_Pos_672 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_672   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_672 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E672_C1_L_Pos and PEAK_C1_Pos <= s_E672_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_672 <= s_Energy_Bin_Pos_672 +'1';
		 Energy_Bin_Pos_Rdy_672 <= '1';
		else
		 s_Energy_Bin_Pos_672 <= s_Energy_Bin_Pos_672;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_672 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_672;   
  
  Energy_Bin_Pos_673 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_673   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_673 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E673_C1_L_Pos and PEAK_C1_Pos <= s_E673_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_673 <= s_Energy_Bin_Pos_673 +'1';
		 Energy_Bin_Pos_Rdy_673 <= '1';
		else
		 s_Energy_Bin_Pos_673 <= s_Energy_Bin_Pos_673;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_673 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_673;   
  
  Energy_Bin_Pos_674 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_674   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_674 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E674_C1_L_Pos and PEAK_C1_Pos <= s_E674_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_674 <= s_Energy_Bin_Pos_674 +'1';
		 Energy_Bin_Pos_Rdy_674 <= '1';
		else
		 s_Energy_Bin_Pos_674 <= s_Energy_Bin_Pos_674;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_674 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_674;   
 
 
  Energy_Bin_Pos_675 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_675   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_675 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E675_C1_L_Pos and PEAK_C1_Pos <= s_E675_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_675 <= s_Energy_Bin_Pos_675 +'1';
		 Energy_Bin_Pos_Rdy_675 <= '1';
		else
		 s_Energy_Bin_Pos_675 <= s_Energy_Bin_Pos_675;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_675 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_675;  
 
  
  Energy_Bin_Pos_676 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_676   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_676 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E676_C1_L_Pos and PEAK_C1_Pos <= s_E676_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_676 <= s_Energy_Bin_Pos_676 +'1';
		 Energy_Bin_Pos_Rdy_676 <= '1';
		else
		 s_Energy_Bin_Pos_676 <= s_Energy_Bin_Pos_676;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_676 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_676;   
  
 Energy_Bin_Pos_677 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_677   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_677 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E677_C1_L_Pos and PEAK_C1_Pos <= s_E677_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_677 <= s_Energy_Bin_Pos_677 +'1';
		 Energy_Bin_Pos_Rdy_677 <= '1';
		else
		 s_Energy_Bin_Pos_677 <= s_Energy_Bin_Pos_677;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_677 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_677;   
  
  Energy_Bin_Pos_678 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_678   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_678 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E678_C1_L_Pos and PEAK_C1_Pos <= s_E678_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_678 <= s_Energy_Bin_Pos_678 +'1';
		 Energy_Bin_Pos_Rdy_678 <= '1';
		else
		 s_Energy_Bin_Pos_678 <= s_Energy_Bin_Pos_678;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_678 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_678;   
  
  Energy_Bin_Pos_679 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_679   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_679 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E679_C1_L_Pos and PEAK_C1_Pos <= s_E679_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_679 <= s_Energy_Bin_Pos_679 +'1';
		 Energy_Bin_Pos_Rdy_679 <= '1';
		else
		 s_Energy_Bin_Pos_679 <= s_Energy_Bin_Pos_679;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_679 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_679;       
  
     Energy_Bin_Pos_680 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_680   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_680 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E680_C1_L_Pos and PEAK_C1_Pos <= s_E680_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_680 <= s_Energy_Bin_Pos_680 +'1';
		 Energy_Bin_Pos_Rdy_680 <= '1';
		else
		 s_Energy_Bin_Pos_680 <= s_Energy_Bin_Pos_680;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_680 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_680;    
  
  Energy_Bin_Pos_681 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_681   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_681 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E681_C1_L_Pos and PEAK_C1_Pos <= s_E681_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_681 <= s_Energy_Bin_Pos_681 +'1';
		 Energy_Bin_Pos_Rdy_681 <= '1';
		else
		 s_Energy_Bin_Pos_681 <= s_Energy_Bin_Pos_681;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_681 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_681;   
  
  Energy_Bin_Pos_682 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_682   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_682 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E682_C1_L_Pos and PEAK_C1_Pos <= s_E682_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_682 <= s_Energy_Bin_Pos_682 +'1';
		 Energy_Bin_Pos_Rdy_682 <= '1';
		else
		 s_Energy_Bin_Pos_682 <= s_Energy_Bin_Pos_682;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_682 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_682;   
  
  Energy_Bin_Pos_683 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_683   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_683 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E683_C1_L_Pos and PEAK_C1_Pos <= s_E683_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_683 <= s_Energy_Bin_Pos_683 +'1';
		 Energy_Bin_Pos_Rdy_683 <= '1';
		else
		 s_Energy_Bin_Pos_683 <= s_Energy_Bin_Pos_683;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_683 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_683;   
  
  Energy_Bin_Pos_684 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_684   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_684 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E684_C1_L_Pos and PEAK_C1_Pos <= s_E684_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_684 <= s_Energy_Bin_Pos_684 +'1';
		 Energy_Bin_Pos_Rdy_684 <= '1';
		else
		 s_Energy_Bin_Pos_684 <= s_Energy_Bin_Pos_684;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_684 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_684;   
 
 
  Energy_Bin_Pos_685 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_685   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_685 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E685_C1_L_Pos and PEAK_C1_Pos <= s_E685_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_685 <= s_Energy_Bin_Pos_685 +'1';
		 Energy_Bin_Pos_Rdy_685 <= '1';
		else
		 s_Energy_Bin_Pos_685 <= s_Energy_Bin_Pos_685;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_685 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_685;  
 
  
  Energy_Bin_Pos_686 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_686   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_686 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E686_C1_L_Pos and PEAK_C1_Pos <= s_E686_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_686 <= s_Energy_Bin_Pos_686 +'1';
		 Energy_Bin_Pos_Rdy_686 <= '1';
		else
		 s_Energy_Bin_Pos_686 <= s_Energy_Bin_Pos_686;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_686 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_686;   
  
 Energy_Bin_Pos_687 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_687   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_687 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E687_C1_L_Pos and PEAK_C1_Pos <= s_E687_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_687 <= s_Energy_Bin_Pos_687 +'1';
		 Energy_Bin_Pos_Rdy_687 <= '1';
		else
		 s_Energy_Bin_Pos_687 <= s_Energy_Bin_Pos_687;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_687 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_687;   
  
  Energy_Bin_Pos_688 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_688   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_688 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E688_C1_L_Pos and PEAK_C1_Pos <= s_E688_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_688 <= s_Energy_Bin_Pos_688 +'1';
		 Energy_Bin_Pos_Rdy_688 <= '1';
		else
		 s_Energy_Bin_Pos_688 <= s_Energy_Bin_Pos_688;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_688 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_688;   
  
  Energy_Bin_Pos_689 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_689   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_689 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E689_C1_L_Pos and PEAK_C1_Pos <= s_E689_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_689 <= s_Energy_Bin_Pos_689 +'1';
		 Energy_Bin_Pos_Rdy_689 <= '1';
		else
		 s_Energy_Bin_Pos_689 <= s_Energy_Bin_Pos_689;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_689 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_689;      
  
     Energy_Bin_Pos_690 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_690   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_690 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E690_C1_L_Pos and PEAK_C1_Pos <= s_E690_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_690 <= s_Energy_Bin_Pos_690 +'1';
		 Energy_Bin_Pos_Rdy_690 <= '1';
		else
		 s_Energy_Bin_Pos_690 <= s_Energy_Bin_Pos_690;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_690 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_690;    
  
  Energy_Bin_Pos_691 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_691   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_691 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E691_C1_L_Pos and PEAK_C1_Pos <= s_E691_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_691 <= s_Energy_Bin_Pos_691 +'1';
		 Energy_Bin_Pos_Rdy_691 <= '1';
		else
		 s_Energy_Bin_Pos_691 <= s_Energy_Bin_Pos_691;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_691 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_691;   
  
  Energy_Bin_Pos_692 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_692   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_692 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E692_C1_L_Pos and PEAK_C1_Pos <= s_E692_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_692 <= s_Energy_Bin_Pos_692 +'1';
		 Energy_Bin_Pos_Rdy_692 <= '1';
		else
		 s_Energy_Bin_Pos_692 <= s_Energy_Bin_Pos_692;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_692 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_692;   
  
  Energy_Bin_Pos_693 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_693   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_693 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E693_C1_L_Pos and PEAK_C1_Pos <= s_E693_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_693 <= s_Energy_Bin_Pos_693 +'1';
		 Energy_Bin_Pos_Rdy_693 <= '1';
		else
		 s_Energy_Bin_Pos_693 <= s_Energy_Bin_Pos_693;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_693 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_693;   
  
  Energy_Bin_Pos_694 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_694   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_694 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E694_C1_L_Pos and PEAK_C1_Pos <= s_E694_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_694 <= s_Energy_Bin_Pos_694 +'1';
		 Energy_Bin_Pos_Rdy_694 <= '1';
		else
		 s_Energy_Bin_Pos_694 <= s_Energy_Bin_Pos_694;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_694 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_694;   
 
 
  Energy_Bin_Pos_695 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_695   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_695 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E695_C1_L_Pos and PEAK_C1_Pos <= s_E695_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_695 <= s_Energy_Bin_Pos_695 +'1';
		 Energy_Bin_Pos_Rdy_695 <= '1';
		else
		 s_Energy_Bin_Pos_695 <= s_Energy_Bin_Pos_695;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_695 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_695;  
 
  
  Energy_Bin_Pos_696 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_696   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_696 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E696_C1_L_Pos and PEAK_C1_Pos <= s_E696_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_696 <= s_Energy_Bin_Pos_696 +'1';
		 Energy_Bin_Pos_Rdy_696 <= '1';
		else
		 s_Energy_Bin_Pos_696 <= s_Energy_Bin_Pos_696;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_696 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_696;   
  
 Energy_Bin_Pos_697 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_697   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_697 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E697_C1_L_Pos and PEAK_C1_Pos <= s_E697_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_697 <= s_Energy_Bin_Pos_697 +'1';
		 Energy_Bin_Pos_Rdy_697 <= '1';
		else
		 s_Energy_Bin_Pos_697 <= s_Energy_Bin_Pos_697;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_697 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_697;   
  
  Energy_Bin_Pos_698 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_698   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_698 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E698_C1_L_Pos and PEAK_C1_Pos <= s_E698_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_698 <= s_Energy_Bin_Pos_698 +'1';
		 Energy_Bin_Pos_Rdy_698 <= '1';
		else
		 s_Energy_Bin_Pos_698 <= s_Energy_Bin_Pos_698;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_698 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_698;   
  
  Energy_Bin_Pos_699 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_699   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_699 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E699_C1_L_Pos and PEAK_C1_Pos <= s_E699_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_699 <= s_Energy_Bin_Pos_699 +'1';
		 Energy_Bin_Pos_Rdy_699 <= '1';
		else
		 s_Energy_Bin_Pos_699 <= s_Energy_Bin_Pos_699;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_699 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_699;   

    Energy_Bin_Pos_700 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_700   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_700 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E700_C1_L_Pos and PEAK_C1_Pos <= s_E700_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_700 <= s_Energy_Bin_Pos_700 +'1';
		 Energy_Bin_Pos_Rdy_700 <= '1';
		else
		 s_Energy_Bin_Pos_700 <= s_Energy_Bin_Pos_700;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_700 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_700;    
  
  Energy_Bin_Pos_701 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_701   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_701 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E701_C1_L_Pos and PEAK_C1_Pos <= s_E701_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_701 <= s_Energy_Bin_Pos_701 +'1';
		 Energy_Bin_Pos_Rdy_701 <= '1';
		else
		 s_Energy_Bin_Pos_701 <= s_Energy_Bin_Pos_701;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_701 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_701;   
  
  Energy_Bin_Pos_702 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_702   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_702 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E702_C1_L_Pos and PEAK_C1_Pos <= s_E702_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_702 <= s_Energy_Bin_Pos_702 +'1';
		 Energy_Bin_Pos_Rdy_702 <= '1';
		else
		 s_Energy_Bin_Pos_702 <= s_Energy_Bin_Pos_702;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_702 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_702;   
  
  Energy_Bin_Pos_703 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_703   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_703 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E703_C1_L_Pos and PEAK_C1_Pos <= s_E703_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_703 <= s_Energy_Bin_Pos_703 +'1';
		 Energy_Bin_Pos_Rdy_703 <= '1';
		else
		 s_Energy_Bin_Pos_703 <= s_Energy_Bin_Pos_703;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_703 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_703;   
  
  Energy_Bin_Pos_704 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_704   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_704 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E704_C1_L_Pos and PEAK_C1_Pos <= s_E704_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_704 <= s_Energy_Bin_Pos_704 +'1';
		 Energy_Bin_Pos_Rdy_704 <= '1';
		else
		 s_Energy_Bin_Pos_704 <= s_Energy_Bin_Pos_704;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_704 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_704;   
 
 
  Energy_Bin_Pos_705 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_705   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_705 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E705_C1_L_Pos and PEAK_C1_Pos <= s_E705_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_705 <= s_Energy_Bin_Pos_705 +'1';
		 Energy_Bin_Pos_Rdy_705 <= '1';
		else
		 s_Energy_Bin_Pos_705 <= s_Energy_Bin_Pos_705;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_705 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_705;  
 
  
  Energy_Bin_Pos_706 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_706   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_706 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E706_C1_L_Pos and PEAK_C1_Pos <= s_E706_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_706 <= s_Energy_Bin_Pos_706 +'1';
		 Energy_Bin_Pos_Rdy_706 <= '1';
		else
		 s_Energy_Bin_Pos_706 <= s_Energy_Bin_Pos_706;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_706 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_706;   
  
 Energy_Bin_Pos_707 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_707   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_707 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E707_C1_L_Pos and PEAK_C1_Pos <= s_E707_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_707 <= s_Energy_Bin_Pos_707 +'1';
		 Energy_Bin_Pos_Rdy_707 <= '1';
		else
		 s_Energy_Bin_Pos_707 <= s_Energy_Bin_Pos_707;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_707 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_707;   
  
  Energy_Bin_Pos_708 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_708   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_708 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E708_C1_L_Pos and PEAK_C1_Pos <= s_E708_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_708 <= s_Energy_Bin_Pos_708 +'1';
		 Energy_Bin_Pos_Rdy_708 <= '1';
		else
		 s_Energy_Bin_Pos_708 <= s_Energy_Bin_Pos_708;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_708 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_708;   
  
  Energy_Bin_Pos_709 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_709   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_709 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E709_C1_L_Pos and PEAK_C1_Pos <= s_E709_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_709 <= s_Energy_Bin_Pos_709 +'1';
		 Energy_Bin_Pos_Rdy_709 <= '1';
		else
		 s_Energy_Bin_Pos_709 <= s_Energy_Bin_Pos_709;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_709 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_709;      
  
     Energy_Bin_Pos_710 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_710   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_710 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E710_C1_L_Pos and PEAK_C1_Pos <= s_E710_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_710 <= s_Energy_Bin_Pos_710 +'1';
		 Energy_Bin_Pos_Rdy_710 <= '1';
		else
		 s_Energy_Bin_Pos_710 <= s_Energy_Bin_Pos_710;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_710 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_710;    
  
  Energy_Bin_Pos_711 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_711   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_711 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E711_C1_L_Pos and PEAK_C1_Pos <= s_E711_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_711 <= s_Energy_Bin_Pos_711 +'1';
		 Energy_Bin_Pos_Rdy_711 <= '1';
		else
		 s_Energy_Bin_Pos_711 <= s_Energy_Bin_Pos_711;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_711 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_711;   
  
  Energy_Bin_Pos_712 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_712   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_712 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E712_C1_L_Pos and PEAK_C1_Pos <= s_E712_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_712 <= s_Energy_Bin_Pos_712 +'1';
		 Energy_Bin_Pos_Rdy_712 <= '1';
		else
		 s_Energy_Bin_Pos_712 <= s_Energy_Bin_Pos_712;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_712 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_712;   
  
  Energy_Bin_Pos_713 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_713   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_713 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E713_C1_L_Pos and PEAK_C1_Pos <= s_E713_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_713 <= s_Energy_Bin_Pos_713 +'1';
		 Energy_Bin_Pos_Rdy_713 <= '1';
		else
		 s_Energy_Bin_Pos_713 <= s_Energy_Bin_Pos_713;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_713 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_713;   
  
  Energy_Bin_Pos_714 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_714   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_714 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E714_C1_L_Pos and PEAK_C1_Pos <= s_E714_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_714 <= s_Energy_Bin_Pos_714 +'1';
		 Energy_Bin_Pos_Rdy_714 <= '1';
		else
		 s_Energy_Bin_Pos_714 <= s_Energy_Bin_Pos_714;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_714 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_714;   
 
 
  Energy_Bin_Pos_715 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_715   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_715 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E715_C1_L_Pos and PEAK_C1_Pos <= s_E715_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_715 <= s_Energy_Bin_Pos_715 +'1';
		 Energy_Bin_Pos_Rdy_715 <= '1';
		else
		 s_Energy_Bin_Pos_715 <= s_Energy_Bin_Pos_715;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_715 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_715;  
 
  
  Energy_Bin_Pos_716 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_716   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_716 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E716_C1_L_Pos and PEAK_C1_Pos <= s_E716_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_716 <= s_Energy_Bin_Pos_716 +'1';
		 Energy_Bin_Pos_Rdy_716 <= '1';
		else
		 s_Energy_Bin_Pos_716 <= s_Energy_Bin_Pos_716;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_716 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_716;   
  
 Energy_Bin_Pos_717 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_717   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_717 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E717_C1_L_Pos and PEAK_C1_Pos <= s_E717_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_717 <= s_Energy_Bin_Pos_717 +'1';
		 Energy_Bin_Pos_Rdy_717 <= '1';
		else
		 s_Energy_Bin_Pos_717 <= s_Energy_Bin_Pos_717;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_717 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_717;   
  
  Energy_Bin_Pos_718 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_718   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_718 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E718_C1_L_Pos and PEAK_C1_Pos <= s_E718_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_718 <= s_Energy_Bin_Pos_718 +'1';
		 Energy_Bin_Pos_Rdy_718 <= '1';
		else
		 s_Energy_Bin_Pos_718 <= s_Energy_Bin_Pos_718;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_718 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_718;   
  
  Energy_Bin_Pos_719 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_719   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_719 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E719_C1_L_Pos and PEAK_C1_Pos <= s_E719_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_719 <= s_Energy_Bin_Pos_719 +'1';
		 Energy_Bin_Pos_Rdy_719 <= '1';
		else
		 s_Energy_Bin_Pos_719 <= s_Energy_Bin_Pos_719;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_719 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_719;       
  
     Energy_Bin_Pos_720 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_720   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_720 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E720_C1_L_Pos and PEAK_C1_Pos <= s_E720_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_720 <= s_Energy_Bin_Pos_720 +'1';
		 Energy_Bin_Pos_Rdy_720 <= '1';
		else
		 s_Energy_Bin_Pos_720 <= s_Energy_Bin_Pos_720;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_720 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_720;    
  
  Energy_Bin_Pos_721 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_721   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_721 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E721_C1_L_Pos and PEAK_C1_Pos <= s_E721_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_721 <= s_Energy_Bin_Pos_721 +'1';
		 Energy_Bin_Pos_Rdy_721 <= '1';
		else
		 s_Energy_Bin_Pos_721 <= s_Energy_Bin_Pos_721;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_721 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_721;   
  
  Energy_Bin_Pos_722 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_722   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_722 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E722_C1_L_Pos and PEAK_C1_Pos <= s_E722_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_722 <= s_Energy_Bin_Pos_722 +'1';
		 Energy_Bin_Pos_Rdy_722 <= '1';
		else
		 s_Energy_Bin_Pos_722 <= s_Energy_Bin_Pos_722;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_722 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_722;   
  
  Energy_Bin_Pos_723 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_723   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_723 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E723_C1_L_Pos and PEAK_C1_Pos <= s_E723_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_723 <= s_Energy_Bin_Pos_723 +'1';
		 Energy_Bin_Pos_Rdy_723 <= '1';
		else
		 s_Energy_Bin_Pos_723 <= s_Energy_Bin_Pos_723;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_723 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_723;   
  
  Energy_Bin_Pos_724 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_724   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_724 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E724_C1_L_Pos and PEAK_C1_Pos <= s_E724_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_724 <= s_Energy_Bin_Pos_724 +'1';
		 Energy_Bin_Pos_Rdy_724 <= '1';
		else
		 s_Energy_Bin_Pos_724 <= s_Energy_Bin_Pos_724;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_724 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_724;   
 
 
  Energy_Bin_Pos_725 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_725   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_725 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E725_C1_L_Pos and PEAK_C1_Pos <= s_E725_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_725 <= s_Energy_Bin_Pos_725 +'1';
		 Energy_Bin_Pos_Rdy_725 <= '1';
		else
		 s_Energy_Bin_Pos_725 <= s_Energy_Bin_Pos_725;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_725 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_725;  
 
  
  Energy_Bin_Pos_726 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_726   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_726 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E726_C1_L_Pos and PEAK_C1_Pos <= s_E726_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_726 <= s_Energy_Bin_Pos_726 +'1';
		 Energy_Bin_Pos_Rdy_726 <= '1';
		else
		 s_Energy_Bin_Pos_726 <= s_Energy_Bin_Pos_726;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_726 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_726;   
  
 Energy_Bin_Pos_727 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_727   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_727 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E727_C1_L_Pos and PEAK_C1_Pos <= s_E727_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_727 <= s_Energy_Bin_Pos_727 +'1';
		 Energy_Bin_Pos_Rdy_727 <= '1';
		else
		 s_Energy_Bin_Pos_727 <= s_Energy_Bin_Pos_727;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_727 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_727;   
  
  Energy_Bin_Pos_728 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_728   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_728 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E728_C1_L_Pos and PEAK_C1_Pos <= s_E728_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_728 <= s_Energy_Bin_Pos_728 +'1';
		 Energy_Bin_Pos_Rdy_728 <= '1';
		else
		 s_Energy_Bin_Pos_728 <= s_Energy_Bin_Pos_728;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_728 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_728;   
  
  Energy_Bin_Pos_729 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_729   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_729 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E729_C1_L_Pos and PEAK_C1_Pos <= s_E729_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_729 <= s_Energy_Bin_Pos_729 +'1';
		 Energy_Bin_Pos_Rdy_729 <= '1';
		else
		 s_Energy_Bin_Pos_729 <= s_Energy_Bin_Pos_729;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_729 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_729;        
  
     Energy_Bin_Pos_730 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_730   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_730 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E730_C1_L_Pos and PEAK_C1_Pos <= s_E730_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_730 <= s_Energy_Bin_Pos_730 +'1';
		 Energy_Bin_Pos_Rdy_730 <= '1';
		else
		 s_Energy_Bin_Pos_730 <= s_Energy_Bin_Pos_730;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_730 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_730;    
  
  Energy_Bin_Pos_731 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_731   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_731 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E731_C1_L_Pos and PEAK_C1_Pos <= s_E731_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_731 <= s_Energy_Bin_Pos_731 +'1';
		 Energy_Bin_Pos_Rdy_731 <= '1';
		else
		 s_Energy_Bin_Pos_731 <= s_Energy_Bin_Pos_731;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_731 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_731;   
  
  Energy_Bin_Pos_732 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_732   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_732 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E732_C1_L_Pos and PEAK_C1_Pos <= s_E732_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_732 <= s_Energy_Bin_Pos_732 +'1';
		 Energy_Bin_Pos_Rdy_732 <= '1';
		else
		 s_Energy_Bin_Pos_732 <= s_Energy_Bin_Pos_732;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_732 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_732;   
  
  Energy_Bin_Pos_733 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_733   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_733 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E733_C1_L_Pos and PEAK_C1_Pos <= s_E733_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_733 <= s_Energy_Bin_Pos_733 +'1';
		 Energy_Bin_Pos_Rdy_733 <= '1';
		else
		 s_Energy_Bin_Pos_733 <= s_Energy_Bin_Pos_733;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_733 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_733;   
  
  Energy_Bin_Pos_734 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_734   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_734 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E734_C1_L_Pos and PEAK_C1_Pos <= s_E734_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_734 <= s_Energy_Bin_Pos_734 +'1';
		 Energy_Bin_Pos_Rdy_734 <= '1';
		else
		 s_Energy_Bin_Pos_734 <= s_Energy_Bin_Pos_734;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_734 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_734;   
 
 
  Energy_Bin_Pos_735 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_735   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_735 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E735_C1_L_Pos and PEAK_C1_Pos <= s_E735_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_735 <= s_Energy_Bin_Pos_735 +'1';
		 Energy_Bin_Pos_Rdy_735 <= '1';
		else
		 s_Energy_Bin_Pos_735 <= s_Energy_Bin_Pos_735;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_735 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_735;  
 
  
  Energy_Bin_Pos_736 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_736   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_736 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E736_C1_L_Pos and PEAK_C1_Pos <= s_E736_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_736 <= s_Energy_Bin_Pos_736 +'1';
		 Energy_Bin_Pos_Rdy_736 <= '1';
		else
		 s_Energy_Bin_Pos_736 <= s_Energy_Bin_Pos_736;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_736 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_736;   
  
 Energy_Bin_Pos_737 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_737   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_737 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E737_C1_L_Pos and PEAK_C1_Pos <= s_E737_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_737 <= s_Energy_Bin_Pos_737 +'1';
		 Energy_Bin_Pos_Rdy_737 <= '1';
		else
		 s_Energy_Bin_Pos_737 <= s_Energy_Bin_Pos_737;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_737 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_737;   
  
  Energy_Bin_Pos_738 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_738   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_738 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E738_C1_L_Pos and PEAK_C1_Pos <= s_E738_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_738 <= s_Energy_Bin_Pos_738 +'1';
		 Energy_Bin_Pos_Rdy_738 <= '1';
		else
		 s_Energy_Bin_Pos_738 <= s_Energy_Bin_Pos_738;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_738 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_738;   
  
  Energy_Bin_Pos_739 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_739   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_739 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E739_C1_L_Pos and PEAK_C1_Pos <= s_E739_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_739 <= s_Energy_Bin_Pos_739 +'1';
		 Energy_Bin_Pos_Rdy_739 <= '1';
		else
		 s_Energy_Bin_Pos_739 <= s_Energy_Bin_Pos_739;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_739 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_739;         
  
     Energy_Bin_Pos_740 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_740   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_740 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E740_C1_L_Pos and PEAK_C1_Pos <= s_E740_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_740 <= s_Energy_Bin_Pos_740 +'1';
		 Energy_Bin_Pos_Rdy_740 <= '1';
		else
		 s_Energy_Bin_Pos_740 <= s_Energy_Bin_Pos_740;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_740 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_740;    
  
  Energy_Bin_Pos_741 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_741   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_741 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E741_C1_L_Pos and PEAK_C1_Pos <= s_E741_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_741 <= s_Energy_Bin_Pos_741 +'1';
		 Energy_Bin_Pos_Rdy_741 <= '1';
		else
		 s_Energy_Bin_Pos_741 <= s_Energy_Bin_Pos_741;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_741 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_741;   
  
  Energy_Bin_Pos_742 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_742   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_742 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E742_C1_L_Pos and PEAK_C1_Pos <= s_E742_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_742 <= s_Energy_Bin_Pos_742 +'1';
		 Energy_Bin_Pos_Rdy_742 <= '1';
		else
		 s_Energy_Bin_Pos_742 <= s_Energy_Bin_Pos_742;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_742 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_742;   
  
  Energy_Bin_Pos_743 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_743   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_743 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E743_C1_L_Pos and PEAK_C1_Pos <= s_E743_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_743 <= s_Energy_Bin_Pos_743 +'1';
		 Energy_Bin_Pos_Rdy_743 <= '1';
		else
		 s_Energy_Bin_Pos_743 <= s_Energy_Bin_Pos_743;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_743 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_743;   
  
  Energy_Bin_Pos_744 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_744   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_744 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E744_C1_L_Pos and PEAK_C1_Pos <= s_E744_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_744 <= s_Energy_Bin_Pos_744 +'1';
		 Energy_Bin_Pos_Rdy_744 <= '1';
		else
		 s_Energy_Bin_Pos_744 <= s_Energy_Bin_Pos_744;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_744 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_744;   
 
 
  Energy_Bin_Pos_745 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_745   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_745 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E745_C1_L_Pos and PEAK_C1_Pos <= s_E745_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_745 <= s_Energy_Bin_Pos_745 +'1';
		 Energy_Bin_Pos_Rdy_745 <= '1';
		else
		 s_Energy_Bin_Pos_745 <= s_Energy_Bin_Pos_745;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_745 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_745;  
 
  
  Energy_Bin_Pos_746 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_746   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_746 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E746_C1_L_Pos and PEAK_C1_Pos <= s_E746_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_746 <= s_Energy_Bin_Pos_746 +'1';
		 Energy_Bin_Pos_Rdy_746 <= '1';
		else
		 s_Energy_Bin_Pos_746 <= s_Energy_Bin_Pos_746;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_746 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_746;   
  
 Energy_Bin_Pos_747 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_747   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_747 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E747_C1_L_Pos and PEAK_C1_Pos <= s_E747_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_747 <= s_Energy_Bin_Pos_747 +'1';
		 Energy_Bin_Pos_Rdy_747 <= '1';
		else
		 s_Energy_Bin_Pos_747 <= s_Energy_Bin_Pos_747;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_747 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_747;   
  
  Energy_Bin_Pos_748 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_748   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_748 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E748_C1_L_Pos and PEAK_C1_Pos <= s_E748_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_748 <= s_Energy_Bin_Pos_748 +'1';
		 Energy_Bin_Pos_Rdy_748 <= '1';
		else
		 s_Energy_Bin_Pos_748 <= s_Energy_Bin_Pos_748;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_748 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_748;   
  
  Energy_Bin_Pos_749 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_749   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_749 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E749_C1_L_Pos and PEAK_C1_Pos <= s_E749_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_749 <= s_Energy_Bin_Pos_749 +'1';
		 Energy_Bin_Pos_Rdy_749 <= '1';
		else
		 s_Energy_Bin_Pos_749 <= s_Energy_Bin_Pos_749;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_749 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_749;          
  
  
     Energy_Bin_Pos_750 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_750   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_750 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E750_C1_L_Pos and PEAK_C1_Pos <= s_E750_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_750 <= s_Energy_Bin_Pos_750 +'1';
		 Energy_Bin_Pos_Rdy_750 <= '1';
		else
		 s_Energy_Bin_Pos_750 <= s_Energy_Bin_Pos_750;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_750 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_750;    
  
  Energy_Bin_Pos_751 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_751   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_751 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E751_C1_L_Pos and PEAK_C1_Pos <= s_E751_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_751 <= s_Energy_Bin_Pos_751 +'1';
		 Energy_Bin_Pos_Rdy_751 <= '1';
		else
		 s_Energy_Bin_Pos_751 <= s_Energy_Bin_Pos_751;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_751 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_751;   
  
  Energy_Bin_Pos_752 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_752   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_752 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E752_C1_L_Pos and PEAK_C1_Pos <= s_E752_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_752 <= s_Energy_Bin_Pos_752 +'1';
		 Energy_Bin_Pos_Rdy_752 <= '1';
		else
		 s_Energy_Bin_Pos_752 <= s_Energy_Bin_Pos_752;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_752 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_752;   
  
  Energy_Bin_Pos_753 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_753   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_753 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E753_C1_L_Pos and PEAK_C1_Pos <= s_E753_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_753 <= s_Energy_Bin_Pos_753 +'1';
		 Energy_Bin_Pos_Rdy_753 <= '1';
		else
		 s_Energy_Bin_Pos_753 <= s_Energy_Bin_Pos_753;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_753 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_753;   
  
  Energy_Bin_Pos_754 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_754   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_754 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E754_C1_L_Pos and PEAK_C1_Pos <= s_E754_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_754 <= s_Energy_Bin_Pos_754 +'1';
		 Energy_Bin_Pos_Rdy_754 <= '1';
		else
		 s_Energy_Bin_Pos_754 <= s_Energy_Bin_Pos_754;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_754 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_754;   
 
 
  Energy_Bin_Pos_755 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_755   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_755 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E755_C1_L_Pos and PEAK_C1_Pos <= s_E755_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_755 <= s_Energy_Bin_Pos_755 +'1';
		 Energy_Bin_Pos_Rdy_755 <= '1';
		else
		 s_Energy_Bin_Pos_755 <= s_Energy_Bin_Pos_755;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_755 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_755;  
 
  
  Energy_Bin_Pos_756 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_756   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_756 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E756_C1_L_Pos and PEAK_C1_Pos <= s_E756_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_756 <= s_Energy_Bin_Pos_756 +'1';
		 Energy_Bin_Pos_Rdy_756 <= '1';
		else
		 s_Energy_Bin_Pos_756 <= s_Energy_Bin_Pos_756;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_756 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_756;   
  
 Energy_Bin_Pos_757 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_757   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_757 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E757_C1_L_Pos and PEAK_C1_Pos <= s_E757_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_757 <= s_Energy_Bin_Pos_757 +'1';
		 Energy_Bin_Pos_Rdy_757 <= '1';
		else
		 s_Energy_Bin_Pos_757 <= s_Energy_Bin_Pos_757;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_757 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_757;   
  
  Energy_Bin_Pos_758 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_758   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_758 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E758_C1_L_Pos and PEAK_C1_Pos <= s_E758_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_758 <= s_Energy_Bin_Pos_758 +'1';
		 Energy_Bin_Pos_Rdy_758 <= '1';
		else
		 s_Energy_Bin_Pos_758 <= s_Energy_Bin_Pos_758;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_758 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_758;   
  
  Energy_Bin_Pos_759 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_759   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_759 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E759_C1_L_Pos and PEAK_C1_Pos <= s_E759_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_759 <= s_Energy_Bin_Pos_759 +'1';
		 Energy_Bin_Pos_Rdy_759 <= '1';
		else
		 s_Energy_Bin_Pos_759 <= s_Energy_Bin_Pos_759;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_759 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_759;           
  
     Energy_Bin_Pos_760 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_760   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_760 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E760_C1_L_Pos and PEAK_C1_Pos <= s_E760_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_760 <= s_Energy_Bin_Pos_760 +'1';
		 Energy_Bin_Pos_Rdy_760 <= '1';
		else
		 s_Energy_Bin_Pos_760 <= s_Energy_Bin_Pos_760;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_760 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_760;    
  
  Energy_Bin_Pos_761 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_761   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_761 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E761_C1_L_Pos and PEAK_C1_Pos <= s_E761_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_761 <= s_Energy_Bin_Pos_761 +'1';
		 Energy_Bin_Pos_Rdy_761 <= '1';
		else
		 s_Energy_Bin_Pos_761 <= s_Energy_Bin_Pos_761;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_761 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_761;   
  
  Energy_Bin_Pos_762 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_762   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_762 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E762_C1_L_Pos and PEAK_C1_Pos <= s_E762_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_762 <= s_Energy_Bin_Pos_762 +'1';
		 Energy_Bin_Pos_Rdy_762 <= '1';
		else
		 s_Energy_Bin_Pos_762 <= s_Energy_Bin_Pos_762;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_762 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_762;   
  
  Energy_Bin_Pos_763 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_763   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_763 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E763_C1_L_Pos and PEAK_C1_Pos <= s_E763_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_763 <= s_Energy_Bin_Pos_763 +'1';
		 Energy_Bin_Pos_Rdy_763 <= '1';
		else
		 s_Energy_Bin_Pos_763 <= s_Energy_Bin_Pos_763;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_763 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_763;   
  
  Energy_Bin_Pos_764 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_764   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_764 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E764_C1_L_Pos and PEAK_C1_Pos <= s_E764_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_764 <= s_Energy_Bin_Pos_764 +'1';
		 Energy_Bin_Pos_Rdy_764 <= '1';
		else
		 s_Energy_Bin_Pos_764 <= s_Energy_Bin_Pos_764;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_764 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_764;   
 
 
  Energy_Bin_Pos_765 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_765   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_765 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E765_C1_L_Pos and PEAK_C1_Pos <= s_E765_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_765 <= s_Energy_Bin_Pos_765 +'1';
		 Energy_Bin_Pos_Rdy_765 <= '1';
		else
		 s_Energy_Bin_Pos_765 <= s_Energy_Bin_Pos_765;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_765 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_765;  
 
  
  Energy_Bin_Pos_766 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_766   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_766 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E766_C1_L_Pos and PEAK_C1_Pos <= s_E766_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_766 <= s_Energy_Bin_Pos_766 +'1';
		 Energy_Bin_Pos_Rdy_766 <= '1';
		else
		 s_Energy_Bin_Pos_766 <= s_Energy_Bin_Pos_766;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_766 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_766;   
  
 Energy_Bin_Pos_767 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_767   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_767 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E767_C1_L_Pos and PEAK_C1_Pos <= s_E767_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_767 <= s_Energy_Bin_Pos_767 +'1';
		 Energy_Bin_Pos_Rdy_767 <= '1';
		else
		 s_Energy_Bin_Pos_767 <= s_Energy_Bin_Pos_767;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_767 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_767;   
  
  Energy_Bin_Pos_768 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_768   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_768 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E768_C1_L_Pos and PEAK_C1_Pos <= s_E768_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_768 <= s_Energy_Bin_Pos_768 +'1';
		 Energy_Bin_Pos_Rdy_768 <= '1';
		else
		 s_Energy_Bin_Pos_768 <= s_Energy_Bin_Pos_768;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_768 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_768;   
  
  Energy_Bin_Pos_769 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_769   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_769 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E769_C1_L_Pos and PEAK_C1_Pos <= s_E769_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_769 <= s_Energy_Bin_Pos_769 +'1';
		 Energy_Bin_Pos_Rdy_769 <= '1';
		else
		 s_Energy_Bin_Pos_769 <= s_Energy_Bin_Pos_769;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_769 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_769;         
  
     Energy_Bin_Pos_770 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_770   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_770 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E770_C1_L_Pos and PEAK_C1_Pos <= s_E770_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_770 <= s_Energy_Bin_Pos_770 +'1';
		 Energy_Bin_Pos_Rdy_770 <= '1';
		else
		 s_Energy_Bin_Pos_770 <= s_Energy_Bin_Pos_770;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_770 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_770;    
  
  Energy_Bin_Pos_771 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_771   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_771 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E771_C1_L_Pos and PEAK_C1_Pos <= s_E771_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_771 <= s_Energy_Bin_Pos_771 +'1';
		 Energy_Bin_Pos_Rdy_771 <= '1';
		else
		 s_Energy_Bin_Pos_771 <= s_Energy_Bin_Pos_771;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_771 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_771;   
  
  Energy_Bin_Pos_772 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_772   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_772 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E772_C1_L_Pos and PEAK_C1_Pos <= s_E772_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_772 <= s_Energy_Bin_Pos_772 +'1';
		 Energy_Bin_Pos_Rdy_772 <= '1';
		else
		 s_Energy_Bin_Pos_772 <= s_Energy_Bin_Pos_772;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_772 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_772;   
  
  Energy_Bin_Pos_773 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_773   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_773 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E773_C1_L_Pos and PEAK_C1_Pos <= s_E773_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_773 <= s_Energy_Bin_Pos_773 +'1';
		 Energy_Bin_Pos_Rdy_773 <= '1';
		else
		 s_Energy_Bin_Pos_773 <= s_Energy_Bin_Pos_773;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_773 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_773;   
  
  Energy_Bin_Pos_774 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_774   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_774 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E774_C1_L_Pos and PEAK_C1_Pos <= s_E774_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_774 <= s_Energy_Bin_Pos_774 +'1';
		 Energy_Bin_Pos_Rdy_774 <= '1';
		else
		 s_Energy_Bin_Pos_774 <= s_Energy_Bin_Pos_774;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_774 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_774;   
 
 
  Energy_Bin_Pos_775 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_775   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_775 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E775_C1_L_Pos and PEAK_C1_Pos <= s_E775_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_775 <= s_Energy_Bin_Pos_775 +'1';
		 Energy_Bin_Pos_Rdy_775 <= '1';
		else
		 s_Energy_Bin_Pos_775 <= s_Energy_Bin_Pos_775;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_775 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_775;  
 
  
  Energy_Bin_Pos_776 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_776   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_776 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E776_C1_L_Pos and PEAK_C1_Pos <= s_E776_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_776 <= s_Energy_Bin_Pos_776 +'1';
		 Energy_Bin_Pos_Rdy_776 <= '1';
		else
		 s_Energy_Bin_Pos_776 <= s_Energy_Bin_Pos_776;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_776 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_776;   
  
 Energy_Bin_Pos_777 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_777   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_777 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E777_C1_L_Pos and PEAK_C1_Pos <= s_E777_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_777 <= s_Energy_Bin_Pos_777 +'1';
		 Energy_Bin_Pos_Rdy_777 <= '1';
		else
		 s_Energy_Bin_Pos_777 <= s_Energy_Bin_Pos_777;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_777 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_777;   
  
  Energy_Bin_Pos_778 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_778   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_778 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E778_C1_L_Pos and PEAK_C1_Pos <= s_E778_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_778 <= s_Energy_Bin_Pos_778 +'1';
		 Energy_Bin_Pos_Rdy_778 <= '1';
		else
		 s_Energy_Bin_Pos_778 <= s_Energy_Bin_Pos_778;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_778 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_778;   
  
  Energy_Bin_Pos_779 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_779   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_779 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E779_C1_L_Pos and PEAK_C1_Pos <= s_E779_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_779 <= s_Energy_Bin_Pos_779 +'1';
		 Energy_Bin_Pos_Rdy_779 <= '1';
		else
		 s_Energy_Bin_Pos_779 <= s_Energy_Bin_Pos_779;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_779 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_779;       
  
     Energy_Bin_Pos_780 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_780   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_780 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E780_C1_L_Pos and PEAK_C1_Pos <= s_E780_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_780 <= s_Energy_Bin_Pos_780 +'1';
		 Energy_Bin_Pos_Rdy_780 <= '1';
		else
		 s_Energy_Bin_Pos_780 <= s_Energy_Bin_Pos_780;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_780 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_780;    
  
  Energy_Bin_Pos_781 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_781   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_781 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E781_C1_L_Pos and PEAK_C1_Pos <= s_E781_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_781 <= s_Energy_Bin_Pos_781 +'1';
		 Energy_Bin_Pos_Rdy_781 <= '1';
		else
		 s_Energy_Bin_Pos_781 <= s_Energy_Bin_Pos_781;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_781 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_781;   
  
  Energy_Bin_Pos_782 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_782   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_782 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E782_C1_L_Pos and PEAK_C1_Pos <= s_E782_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_782 <= s_Energy_Bin_Pos_782 +'1';
		 Energy_Bin_Pos_Rdy_782 <= '1';
		else
		 s_Energy_Bin_Pos_782 <= s_Energy_Bin_Pos_782;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_782 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_782;   
  
  Energy_Bin_Pos_783 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_783   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_783 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E783_C1_L_Pos and PEAK_C1_Pos <= s_E783_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_783 <= s_Energy_Bin_Pos_783 +'1';
		 Energy_Bin_Pos_Rdy_783 <= '1';
		else
		 s_Energy_Bin_Pos_783 <= s_Energy_Bin_Pos_783;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_783 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_783;   
  
  Energy_Bin_Pos_784 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_784   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_784 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E784_C1_L_Pos and PEAK_C1_Pos <= s_E784_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_784 <= s_Energy_Bin_Pos_784 +'1';
		 Energy_Bin_Pos_Rdy_784 <= '1';
		else
		 s_Energy_Bin_Pos_784 <= s_Energy_Bin_Pos_784;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_784 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_784;   
 
 
  Energy_Bin_Pos_785 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_785   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_785 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E785_C1_L_Pos and PEAK_C1_Pos <= s_E785_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_785 <= s_Energy_Bin_Pos_785 +'1';
		 Energy_Bin_Pos_Rdy_785 <= '1';
		else
		 s_Energy_Bin_Pos_785 <= s_Energy_Bin_Pos_785;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_785 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_785;  
 
  
  Energy_Bin_Pos_786 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_786   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_786 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E786_C1_L_Pos and PEAK_C1_Pos <= s_E786_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_786 <= s_Energy_Bin_Pos_786 +'1';
		 Energy_Bin_Pos_Rdy_786 <= '1';
		else
		 s_Energy_Bin_Pos_786 <= s_Energy_Bin_Pos_786;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_786 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_786;   
  
 Energy_Bin_Pos_787 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_787   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_787 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E787_C1_L_Pos and PEAK_C1_Pos <= s_E787_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_787 <= s_Energy_Bin_Pos_787 +'1';
		 Energy_Bin_Pos_Rdy_787 <= '1';
		else
		 s_Energy_Bin_Pos_787 <= s_Energy_Bin_Pos_787;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_787 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_787;   
  
  Energy_Bin_Pos_788 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_788   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_788 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E788_C1_L_Pos and PEAK_C1_Pos <= s_E788_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_788 <= s_Energy_Bin_Pos_788 +'1';
		 Energy_Bin_Pos_Rdy_788 <= '1';
		else
		 s_Energy_Bin_Pos_788 <= s_Energy_Bin_Pos_788;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_788 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_788;   
  
  Energy_Bin_Pos_789 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_789   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_789 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E789_C1_L_Pos and PEAK_C1_Pos <= s_E789_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_789 <= s_Energy_Bin_Pos_789 +'1';
		 Energy_Bin_Pos_Rdy_789 <= '1';
		else
		 s_Energy_Bin_Pos_789 <= s_Energy_Bin_Pos_789;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_789 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_789;      
  
     Energy_Bin_Pos_790 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_790   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_790 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E790_C1_L_Pos and PEAK_C1_Pos <= s_E790_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_790 <= s_Energy_Bin_Pos_790 +'1';
		 Energy_Bin_Pos_Rdy_790 <= '1';
		else
		 s_Energy_Bin_Pos_790 <= s_Energy_Bin_Pos_790;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_790 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_790;    
  
  Energy_Bin_Pos_791 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_791   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_791 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E791_C1_L_Pos and PEAK_C1_Pos <= s_E791_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_791 <= s_Energy_Bin_Pos_791 +'1';
		 Energy_Bin_Pos_Rdy_791 <= '1';
		else
		 s_Energy_Bin_Pos_791 <= s_Energy_Bin_Pos_791;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_791 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_791;   
  
  Energy_Bin_Pos_792 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_792   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_792 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E792_C1_L_Pos and PEAK_C1_Pos <= s_E792_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_792 <= s_Energy_Bin_Pos_792 +'1';
		 Energy_Bin_Pos_Rdy_792 <= '1';
		else
		 s_Energy_Bin_Pos_792 <= s_Energy_Bin_Pos_792;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_792 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_792;   
  
  Energy_Bin_Pos_793 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_793   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_793 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E793_C1_L_Pos and PEAK_C1_Pos <= s_E793_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_793 <= s_Energy_Bin_Pos_793 +'1';
		 Energy_Bin_Pos_Rdy_793 <= '1';
		else
		 s_Energy_Bin_Pos_793 <= s_Energy_Bin_Pos_793;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_793 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_793;   
  
  Energy_Bin_Pos_794 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_794   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_794 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E794_C1_L_Pos and PEAK_C1_Pos <= s_E794_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_794 <= s_Energy_Bin_Pos_794 +'1';
		 Energy_Bin_Pos_Rdy_794 <= '1';
		else
		 s_Energy_Bin_Pos_794 <= s_Energy_Bin_Pos_794;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_794 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_794;   
 
 
  Energy_Bin_Pos_795 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_795   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_795 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E795_C1_L_Pos and PEAK_C1_Pos <= s_E795_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_795 <= s_Energy_Bin_Pos_795 +'1';
		 Energy_Bin_Pos_Rdy_795 <= '1';
		else
		 s_Energy_Bin_Pos_795 <= s_Energy_Bin_Pos_795;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_795 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_795;  
 
  
  Energy_Bin_Pos_796 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_796   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_796 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E796_C1_L_Pos and PEAK_C1_Pos <= s_E796_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_796 <= s_Energy_Bin_Pos_796 +'1';
		 Energy_Bin_Pos_Rdy_796 <= '1';
		else
		 s_Energy_Bin_Pos_796 <= s_Energy_Bin_Pos_796;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_796 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_796;   
  
 Energy_Bin_Pos_797 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_797   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_797 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E797_C1_L_Pos and PEAK_C1_Pos <= s_E797_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_797 <= s_Energy_Bin_Pos_797 +'1';
		 Energy_Bin_Pos_Rdy_797 <= '1';
		else
		 s_Energy_Bin_Pos_797 <= s_Energy_Bin_Pos_797;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_797 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_797;   
  
  Energy_Bin_Pos_798 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_798   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_798 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E798_C1_L_Pos and PEAK_C1_Pos <= s_E798_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_798 <= s_Energy_Bin_Pos_798 +'1';
		 Energy_Bin_Pos_Rdy_798 <= '1';
		else
		 s_Energy_Bin_Pos_798 <= s_Energy_Bin_Pos_798;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_798 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_798;   
  
  Energy_Bin_Pos_799 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_799   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_799 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E799_C1_L_Pos and PEAK_C1_Pos <= s_E799_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_799 <= s_Energy_Bin_Pos_799 +'1';
		 Energy_Bin_Pos_Rdy_799 <= '1';
		else
		 s_Energy_Bin_Pos_799 <= s_Energy_Bin_Pos_799;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_799 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_799;   

    Energy_Bin_Pos_800 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_800   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_800 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E800_C1_L_Pos and PEAK_C1_Pos <= s_E800_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_800 <= s_Energy_Bin_Pos_800 +'1';
		 Energy_Bin_Pos_Rdy_800 <= '1';
		else
		 s_Energy_Bin_Pos_800 <= s_Energy_Bin_Pos_800;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_800 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_800;    
  
  Energy_Bin_Pos_801 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_801   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_801 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E801_C1_L_Pos and PEAK_C1_Pos <= s_E801_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_801 <= s_Energy_Bin_Pos_801 +'1';
		 Energy_Bin_Pos_Rdy_801 <= '1';
		else
		 s_Energy_Bin_Pos_801 <= s_Energy_Bin_Pos_801;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_801 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_801;   
  
  Energy_Bin_Pos_802 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_802   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_802 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E802_C1_L_Pos and PEAK_C1_Pos <= s_E802_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_802 <= s_Energy_Bin_Pos_802 +'1';
		 Energy_Bin_Pos_Rdy_802 <= '1';
		else
		 s_Energy_Bin_Pos_802 <= s_Energy_Bin_Pos_802;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_802 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_802;   
  
  Energy_Bin_Pos_803 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_803   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_803 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E803_C1_L_Pos and PEAK_C1_Pos <= s_E803_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_803 <= s_Energy_Bin_Pos_803 +'1';
		 Energy_Bin_Pos_Rdy_803 <= '1';
		else
		 s_Energy_Bin_Pos_803 <= s_Energy_Bin_Pos_803;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_803 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_803;   
  
  Energy_Bin_Pos_804 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_804   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_804 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E804_C1_L_Pos and PEAK_C1_Pos <= s_E804_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_804 <= s_Energy_Bin_Pos_804 +'1';
		 Energy_Bin_Pos_Rdy_804 <= '1';
		else
		 s_Energy_Bin_Pos_804 <= s_Energy_Bin_Pos_804;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_804 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_804;   
 
 
  Energy_Bin_Pos_805 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_805   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_805 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E805_C1_L_Pos and PEAK_C1_Pos <= s_E805_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_805 <= s_Energy_Bin_Pos_805 +'1';
		 Energy_Bin_Pos_Rdy_805 <= '1';
		else
		 s_Energy_Bin_Pos_805 <= s_Energy_Bin_Pos_805;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_805 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_805;  
 
  
  Energy_Bin_Pos_806 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_806   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_806 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E806_C1_L_Pos and PEAK_C1_Pos <= s_E806_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_806 <= s_Energy_Bin_Pos_806 +'1';
		 Energy_Bin_Pos_Rdy_806 <= '1';
		else
		 s_Energy_Bin_Pos_806 <= s_Energy_Bin_Pos_806;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_806 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_806;   
  
 Energy_Bin_Pos_807 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_807   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_807 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E807_C1_L_Pos and PEAK_C1_Pos <= s_E807_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_807 <= s_Energy_Bin_Pos_807 +'1';
		 Energy_Bin_Pos_Rdy_807 <= '1';
		else
		 s_Energy_Bin_Pos_807 <= s_Energy_Bin_Pos_807;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_807 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_807;   
  
  Energy_Bin_Pos_808 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_808   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_808 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E808_C1_L_Pos and PEAK_C1_Pos <= s_E808_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_808 <= s_Energy_Bin_Pos_808 +'1';
		 Energy_Bin_Pos_Rdy_808 <= '1';
		else
		 s_Energy_Bin_Pos_808 <= s_Energy_Bin_Pos_808;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_808 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_808;   
  
  Energy_Bin_Pos_809 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_809   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_809 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E809_C1_L_Pos and PEAK_C1_Pos <= s_E809_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_809 <= s_Energy_Bin_Pos_809 +'1';
		 Energy_Bin_Pos_Rdy_809 <= '1';
		else
		 s_Energy_Bin_Pos_809 <= s_Energy_Bin_Pos_809;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_809 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_809;      
  
     Energy_Bin_Pos_810 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_810   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_810 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E810_C1_L_Pos and PEAK_C1_Pos <= s_E810_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_810 <= s_Energy_Bin_Pos_810 +'1';
		 Energy_Bin_Pos_Rdy_810 <= '1';
		else
		 s_Energy_Bin_Pos_810 <= s_Energy_Bin_Pos_810;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_810 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_810;    
  
  Energy_Bin_Pos_811 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_811   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_811 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E811_C1_L_Pos and PEAK_C1_Pos <= s_E811_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_811 <= s_Energy_Bin_Pos_811 +'1';
		 Energy_Bin_Pos_Rdy_811 <= '1';
		else
		 s_Energy_Bin_Pos_811 <= s_Energy_Bin_Pos_811;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_811 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_811;   
  
  Energy_Bin_Pos_812 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_812   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_812 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E812_C1_L_Pos and PEAK_C1_Pos <= s_E812_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_812 <= s_Energy_Bin_Pos_812 +'1';
		 Energy_Bin_Pos_Rdy_812 <= '1';
		else
		 s_Energy_Bin_Pos_812 <= s_Energy_Bin_Pos_812;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_812 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_812;   
  
  Energy_Bin_Pos_813 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_813   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_813 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E813_C1_L_Pos and PEAK_C1_Pos <= s_E813_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_813 <= s_Energy_Bin_Pos_813 +'1';
		 Energy_Bin_Pos_Rdy_813 <= '1';
		else
		 s_Energy_Bin_Pos_813 <= s_Energy_Bin_Pos_813;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_813 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_813;   
  
  Energy_Bin_Pos_814 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_814   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_814 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E814_C1_L_Pos and PEAK_C1_Pos <= s_E814_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_814 <= s_Energy_Bin_Pos_814 +'1';
		 Energy_Bin_Pos_Rdy_814 <= '1';
		else
		 s_Energy_Bin_Pos_814 <= s_Energy_Bin_Pos_814;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_814 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_814;   
 
 
  Energy_Bin_Pos_815 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_815   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_815 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E815_C1_L_Pos and PEAK_C1_Pos <= s_E815_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_815 <= s_Energy_Bin_Pos_815 +'1';
		 Energy_Bin_Pos_Rdy_815 <= '1';
		else
		 s_Energy_Bin_Pos_815 <= s_Energy_Bin_Pos_815;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_815 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_815;  
 
  
  Energy_Bin_Pos_816 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_816   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_816 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E816_C1_L_Pos and PEAK_C1_Pos <= s_E816_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_816 <= s_Energy_Bin_Pos_816 +'1';
		 Energy_Bin_Pos_Rdy_816 <= '1';
		else
		 s_Energy_Bin_Pos_816 <= s_Energy_Bin_Pos_816;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_816 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_816;   
  
 Energy_Bin_Pos_817 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_817   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_817 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E817_C1_L_Pos and PEAK_C1_Pos <= s_E817_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_817 <= s_Energy_Bin_Pos_817 +'1';
		 Energy_Bin_Pos_Rdy_817 <= '1';
		else
		 s_Energy_Bin_Pos_817 <= s_Energy_Bin_Pos_817;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_817 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_817;   
  
  Energy_Bin_Pos_818 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_818   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_818 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E818_C1_L_Pos and PEAK_C1_Pos <= s_E818_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_818 <= s_Energy_Bin_Pos_818 +'1';
		 Energy_Bin_Pos_Rdy_818 <= '1';
		else
		 s_Energy_Bin_Pos_818 <= s_Energy_Bin_Pos_818;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_818 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_818;   
  
  Energy_Bin_Pos_819 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_819   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_819 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E819_C1_L_Pos and PEAK_C1_Pos <= s_E819_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_819 <= s_Energy_Bin_Pos_819 +'1';
		 Energy_Bin_Pos_Rdy_819 <= '1';
		else
		 s_Energy_Bin_Pos_819 <= s_Energy_Bin_Pos_819;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_819 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_819;       
  
     Energy_Bin_Pos_820 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_820   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_820 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E820_C1_L_Pos and PEAK_C1_Pos <= s_E820_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_820 <= s_Energy_Bin_Pos_820 +'1';
		 Energy_Bin_Pos_Rdy_820 <= '1';
		else
		 s_Energy_Bin_Pos_820 <= s_Energy_Bin_Pos_820;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_820 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_820;    
  
  Energy_Bin_Pos_821 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_821   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_821 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E821_C1_L_Pos and PEAK_C1_Pos <= s_E821_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_821 <= s_Energy_Bin_Pos_821 +'1';
		 Energy_Bin_Pos_Rdy_821 <= '1';
		else
		 s_Energy_Bin_Pos_821 <= s_Energy_Bin_Pos_821;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_821 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_821;   
  
  Energy_Bin_Pos_822 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_822   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_822 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E822_C1_L_Pos and PEAK_C1_Pos <= s_E822_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_822 <= s_Energy_Bin_Pos_822 +'1';
		 Energy_Bin_Pos_Rdy_822 <= '1';
		else
		 s_Energy_Bin_Pos_822 <= s_Energy_Bin_Pos_822;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_822 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_822;   
  
  Energy_Bin_Pos_823 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_823   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_823 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E823_C1_L_Pos and PEAK_C1_Pos <= s_E823_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_823 <= s_Energy_Bin_Pos_823 +'1';
		 Energy_Bin_Pos_Rdy_823 <= '1';
		else
		 s_Energy_Bin_Pos_823 <= s_Energy_Bin_Pos_823;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_823 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_823;   
  
  Energy_Bin_Pos_824 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_824   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_824 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E824_C1_L_Pos and PEAK_C1_Pos <= s_E824_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_824 <= s_Energy_Bin_Pos_824 +'1';
		 Energy_Bin_Pos_Rdy_824 <= '1';
		else
		 s_Energy_Bin_Pos_824 <= s_Energy_Bin_Pos_824;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_824 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_824;   
 
 
  Energy_Bin_Pos_825 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_825   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_825 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E825_C1_L_Pos and PEAK_C1_Pos <= s_E825_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_825 <= s_Energy_Bin_Pos_825 +'1';
		 Energy_Bin_Pos_Rdy_825 <= '1';
		else
		 s_Energy_Bin_Pos_825 <= s_Energy_Bin_Pos_825;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_825 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_825;  
 
  
  Energy_Bin_Pos_826 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_826   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_826 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E826_C1_L_Pos and PEAK_C1_Pos <= s_E826_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_826 <= s_Energy_Bin_Pos_826 +'1';
		 Energy_Bin_Pos_Rdy_826 <= '1';
		else
		 s_Energy_Bin_Pos_826 <= s_Energy_Bin_Pos_826;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_826 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_826;   
  
 Energy_Bin_Pos_827 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_827   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_827 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E827_C1_L_Pos and PEAK_C1_Pos <= s_E827_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_827 <= s_Energy_Bin_Pos_827 +'1';
		 Energy_Bin_Pos_Rdy_827 <= '1';
		else
		 s_Energy_Bin_Pos_827 <= s_Energy_Bin_Pos_827;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_827 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_827;   
  
  Energy_Bin_Pos_828 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_828   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_828 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E828_C1_L_Pos and PEAK_C1_Pos <= s_E828_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_828 <= s_Energy_Bin_Pos_828 +'1';
		 Energy_Bin_Pos_Rdy_828 <= '1';
		else
		 s_Energy_Bin_Pos_828 <= s_Energy_Bin_Pos_828;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_828 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_828;   
  
  Energy_Bin_Pos_829 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_829   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_829 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E829_C1_L_Pos and PEAK_C1_Pos <= s_E829_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_829 <= s_Energy_Bin_Pos_829 +'1';
		 Energy_Bin_Pos_Rdy_829 <= '1';
		else
		 s_Energy_Bin_Pos_829 <= s_Energy_Bin_Pos_829;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_829 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_829;        
  
     Energy_Bin_Pos_830 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_830   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_830 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E830_C1_L_Pos and PEAK_C1_Pos <= s_E830_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_830 <= s_Energy_Bin_Pos_830 +'1';
		 Energy_Bin_Pos_Rdy_830 <= '1';
		else
		 s_Energy_Bin_Pos_830 <= s_Energy_Bin_Pos_830;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_830 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_830;    
  
  Energy_Bin_Pos_831 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_831   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_831 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E831_C1_L_Pos and PEAK_C1_Pos <= s_E831_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_831 <= s_Energy_Bin_Pos_831 +'1';
		 Energy_Bin_Pos_Rdy_831 <= '1';
		else
		 s_Energy_Bin_Pos_831 <= s_Energy_Bin_Pos_831;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_831 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_831;   
  
  Energy_Bin_Pos_832 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_832   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_832 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E832_C1_L_Pos and PEAK_C1_Pos <= s_E832_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_832 <= s_Energy_Bin_Pos_832 +'1';
		 Energy_Bin_Pos_Rdy_832 <= '1';
		else
		 s_Energy_Bin_Pos_832 <= s_Energy_Bin_Pos_832;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_832 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_832;   
  
  Energy_Bin_Pos_833 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_833   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_833 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E833_C1_L_Pos and PEAK_C1_Pos <= s_E833_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_833 <= s_Energy_Bin_Pos_833 +'1';
		 Energy_Bin_Pos_Rdy_833 <= '1';
		else
		 s_Energy_Bin_Pos_833 <= s_Energy_Bin_Pos_833;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_833 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_833;   
  
  Energy_Bin_Pos_834 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_834   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_834 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E834_C1_L_Pos and PEAK_C1_Pos <= s_E834_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_834 <= s_Energy_Bin_Pos_834 +'1';
		 Energy_Bin_Pos_Rdy_834 <= '1';
		else
		 s_Energy_Bin_Pos_834 <= s_Energy_Bin_Pos_834;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_834 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_834;   
 
 
  Energy_Bin_Pos_835 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_835   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_835 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E835_C1_L_Pos and PEAK_C1_Pos <= s_E835_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_835 <= s_Energy_Bin_Pos_835 +'1';
		 Energy_Bin_Pos_Rdy_835 <= '1';
		else
		 s_Energy_Bin_Pos_835 <= s_Energy_Bin_Pos_835;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_835 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_835;  
 
  
  Energy_Bin_Pos_836 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_836   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_836 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E836_C1_L_Pos and PEAK_C1_Pos <= s_E836_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_836 <= s_Energy_Bin_Pos_836 +'1';
		 Energy_Bin_Pos_Rdy_836 <= '1';
		else
		 s_Energy_Bin_Pos_836 <= s_Energy_Bin_Pos_836;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_836 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_836;   
  
 Energy_Bin_Pos_837 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_837   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_837 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E837_C1_L_Pos and PEAK_C1_Pos <= s_E837_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_837 <= s_Energy_Bin_Pos_837 +'1';
		 Energy_Bin_Pos_Rdy_837 <= '1';
		else
		 s_Energy_Bin_Pos_837 <= s_Energy_Bin_Pos_837;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_837 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_837;   
  
  Energy_Bin_Pos_838 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_838   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_838 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E838_C1_L_Pos and PEAK_C1_Pos <= s_E838_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_838 <= s_Energy_Bin_Pos_838 +'1';
		 Energy_Bin_Pos_Rdy_838 <= '1';
		else
		 s_Energy_Bin_Pos_838 <= s_Energy_Bin_Pos_838;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_838 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_838;   
  
  Energy_Bin_Pos_839 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_839   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_839 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E839_C1_L_Pos and PEAK_C1_Pos <= s_E839_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_839 <= s_Energy_Bin_Pos_839 +'1';
		 Energy_Bin_Pos_Rdy_839 <= '1';
		else
		 s_Energy_Bin_Pos_839 <= s_Energy_Bin_Pos_839;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_839 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_839;         
  
     Energy_Bin_Pos_840 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_840   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_840 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E840_C1_L_Pos and PEAK_C1_Pos <= s_E840_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_840 <= s_Energy_Bin_Pos_840 +'1';
		 Energy_Bin_Pos_Rdy_840 <= '1';
		else
		 s_Energy_Bin_Pos_840 <= s_Energy_Bin_Pos_840;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_840 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_840;    
  
  Energy_Bin_Pos_841 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_841   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_841 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E841_C1_L_Pos and PEAK_C1_Pos <= s_E841_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_841 <= s_Energy_Bin_Pos_841 +'1';
		 Energy_Bin_Pos_Rdy_841 <= '1';
		else
		 s_Energy_Bin_Pos_841 <= s_Energy_Bin_Pos_841;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_841 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_841;   
  
  Energy_Bin_Pos_842 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_842   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_842 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E842_C1_L_Pos and PEAK_C1_Pos <= s_E842_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_842 <= s_Energy_Bin_Pos_842 +'1';
		 Energy_Bin_Pos_Rdy_842 <= '1';
		else
		 s_Energy_Bin_Pos_842 <= s_Energy_Bin_Pos_842;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_842 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_842;   
  
  Energy_Bin_Pos_843 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_843   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_843 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E843_C1_L_Pos and PEAK_C1_Pos <= s_E843_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_843 <= s_Energy_Bin_Pos_843 +'1';
		 Energy_Bin_Pos_Rdy_843 <= '1';
		else
		 s_Energy_Bin_Pos_843 <= s_Energy_Bin_Pos_843;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_843 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_843;   
  
  Energy_Bin_Pos_844 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_844   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_844 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E844_C1_L_Pos and PEAK_C1_Pos <= s_E844_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_844 <= s_Energy_Bin_Pos_844 +'1';
		 Energy_Bin_Pos_Rdy_844 <= '1';
		else
		 s_Energy_Bin_Pos_844 <= s_Energy_Bin_Pos_844;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_844 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_844;   
 
 
  Energy_Bin_Pos_845 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_845   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_845 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E845_C1_L_Pos and PEAK_C1_Pos <= s_E845_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_845 <= s_Energy_Bin_Pos_845 +'1';
		 Energy_Bin_Pos_Rdy_845 <= '1';
		else
		 s_Energy_Bin_Pos_845 <= s_Energy_Bin_Pos_845;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_845 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_845;  
 
  
  Energy_Bin_Pos_846 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_846   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_846 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E846_C1_L_Pos and PEAK_C1_Pos <= s_E846_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_846 <= s_Energy_Bin_Pos_846 +'1';
		 Energy_Bin_Pos_Rdy_846 <= '1';
		else
		 s_Energy_Bin_Pos_846 <= s_Energy_Bin_Pos_846;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_846 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_846;   
  
 Energy_Bin_Pos_847 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_847   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_847 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E847_C1_L_Pos and PEAK_C1_Pos <= s_E847_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_847 <= s_Energy_Bin_Pos_847 +'1';
		 Energy_Bin_Pos_Rdy_847 <= '1';
		else
		 s_Energy_Bin_Pos_847 <= s_Energy_Bin_Pos_847;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_847 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_847;   
  
  Energy_Bin_Pos_848 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_848   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_848 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E848_C1_L_Pos and PEAK_C1_Pos <= s_E848_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_848 <= s_Energy_Bin_Pos_848 +'1';
		 Energy_Bin_Pos_Rdy_848 <= '1';
		else
		 s_Energy_Bin_Pos_848 <= s_Energy_Bin_Pos_848;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_848 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_848;   
  
  Energy_Bin_Pos_849 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_849   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_849 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E849_C1_L_Pos and PEAK_C1_Pos <= s_E849_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_849 <= s_Energy_Bin_Pos_849 +'1';
		 Energy_Bin_Pos_Rdy_849 <= '1';
		else
		 s_Energy_Bin_Pos_849 <= s_Energy_Bin_Pos_849;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_849 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_849;          
  
  
     Energy_Bin_Pos_850 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_850   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_850 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E850_C1_L_Pos and PEAK_C1_Pos <= s_E850_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_850 <= s_Energy_Bin_Pos_850 +'1';
		 Energy_Bin_Pos_Rdy_850 <= '1';
		else
		 s_Energy_Bin_Pos_850 <= s_Energy_Bin_Pos_850;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_850 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_850;    
  
  Energy_Bin_Pos_851 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_851   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_851 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E851_C1_L_Pos and PEAK_C1_Pos <= s_E851_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_851 <= s_Energy_Bin_Pos_851 +'1';
		 Energy_Bin_Pos_Rdy_851 <= '1';
		else
		 s_Energy_Bin_Pos_851 <= s_Energy_Bin_Pos_851;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_851 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_851;   
  
  Energy_Bin_Pos_852 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_852   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_852 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E852_C1_L_Pos and PEAK_C1_Pos <= s_E852_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_852 <= s_Energy_Bin_Pos_852 +'1';
		 Energy_Bin_Pos_Rdy_852 <= '1';
		else
		 s_Energy_Bin_Pos_852 <= s_Energy_Bin_Pos_852;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_852 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_852;   
  
  Energy_Bin_Pos_853 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_853   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_853 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E853_C1_L_Pos and PEAK_C1_Pos <= s_E853_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_853 <= s_Energy_Bin_Pos_853 +'1';
		 Energy_Bin_Pos_Rdy_853 <= '1';
		else
		 s_Energy_Bin_Pos_853 <= s_Energy_Bin_Pos_853;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_853 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_853;   
  
  Energy_Bin_Pos_854 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_854   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_854 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E854_C1_L_Pos and PEAK_C1_Pos <= s_E854_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_854 <= s_Energy_Bin_Pos_854 +'1';
		 Energy_Bin_Pos_Rdy_854 <= '1';
		else
		 s_Energy_Bin_Pos_854 <= s_Energy_Bin_Pos_854;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_854 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_854;   
 
 
  Energy_Bin_Pos_855 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_855   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_855 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E855_C1_L_Pos and PEAK_C1_Pos <= s_E855_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_855 <= s_Energy_Bin_Pos_855 +'1';
		 Energy_Bin_Pos_Rdy_855 <= '1';
		else
		 s_Energy_Bin_Pos_855 <= s_Energy_Bin_Pos_855;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_855 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_855;  
 
  
  Energy_Bin_Pos_856 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_856   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_856 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E856_C1_L_Pos and PEAK_C1_Pos <= s_E856_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_856 <= s_Energy_Bin_Pos_856 +'1';
		 Energy_Bin_Pos_Rdy_856 <= '1';
		else
		 s_Energy_Bin_Pos_856 <= s_Energy_Bin_Pos_856;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_856 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_856;   
  
 Energy_Bin_Pos_857 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_857   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_857 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E857_C1_L_Pos and PEAK_C1_Pos <= s_E857_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_857 <= s_Energy_Bin_Pos_857 +'1';
		 Energy_Bin_Pos_Rdy_857 <= '1';
		else
		 s_Energy_Bin_Pos_857 <= s_Energy_Bin_Pos_857;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_857 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_857;   
  
  Energy_Bin_Pos_858 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_858   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_858 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E858_C1_L_Pos and PEAK_C1_Pos <= s_E858_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_858 <= s_Energy_Bin_Pos_858 +'1';
		 Energy_Bin_Pos_Rdy_858 <= '1';
		else
		 s_Energy_Bin_Pos_858 <= s_Energy_Bin_Pos_858;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_858 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_858;   
  
  Energy_Bin_Pos_859 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_859   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_859 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E859_C1_L_Pos and PEAK_C1_Pos <= s_E859_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_859 <= s_Energy_Bin_Pos_859 +'1';
		 Energy_Bin_Pos_Rdy_859 <= '1';
		else
		 s_Energy_Bin_Pos_859 <= s_Energy_Bin_Pos_859;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_859 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_859;           
  
     Energy_Bin_Pos_860 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_860   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_860 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E860_C1_L_Pos and PEAK_C1_Pos <= s_E860_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_860 <= s_Energy_Bin_Pos_860 +'1';
		 Energy_Bin_Pos_Rdy_860 <= '1';
		else
		 s_Energy_Bin_Pos_860 <= s_Energy_Bin_Pos_860;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_860 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_860;    
  
  Energy_Bin_Pos_861 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_861   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_861 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E861_C1_L_Pos and PEAK_C1_Pos <= s_E861_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_861 <= s_Energy_Bin_Pos_861 +'1';
		 Energy_Bin_Pos_Rdy_861 <= '1';
		else
		 s_Energy_Bin_Pos_861 <= s_Energy_Bin_Pos_861;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_861 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_861;   
  
  Energy_Bin_Pos_862 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_862   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_862 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E862_C1_L_Pos and PEAK_C1_Pos <= s_E862_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_862 <= s_Energy_Bin_Pos_862 +'1';
		 Energy_Bin_Pos_Rdy_862 <= '1';
		else
		 s_Energy_Bin_Pos_862 <= s_Energy_Bin_Pos_862;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_862 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_862;   
  
  Energy_Bin_Pos_863 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_863   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_863 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E863_C1_L_Pos and PEAK_C1_Pos <= s_E863_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_863 <= s_Energy_Bin_Pos_863 +'1';
		 Energy_Bin_Pos_Rdy_863 <= '1';
		else
		 s_Energy_Bin_Pos_863 <= s_Energy_Bin_Pos_863;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_863 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_863;   
  
  Energy_Bin_Pos_864 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_864   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_864 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E864_C1_L_Pos and PEAK_C1_Pos <= s_E864_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_864 <= s_Energy_Bin_Pos_864 +'1';
		 Energy_Bin_Pos_Rdy_864 <= '1';
		else
		 s_Energy_Bin_Pos_864 <= s_Energy_Bin_Pos_864;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_864 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_864;   
 
 
  Energy_Bin_Pos_865 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_865   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_865 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E865_C1_L_Pos and PEAK_C1_Pos <= s_E865_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_865 <= s_Energy_Bin_Pos_865 +'1';
		 Energy_Bin_Pos_Rdy_865 <= '1';
		else
		 s_Energy_Bin_Pos_865 <= s_Energy_Bin_Pos_865;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_865 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_865;  
 
  
  Energy_Bin_Pos_866 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_866   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_866 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E866_C1_L_Pos and PEAK_C1_Pos <= s_E866_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_866 <= s_Energy_Bin_Pos_866 +'1';
		 Energy_Bin_Pos_Rdy_866 <= '1';
		else
		 s_Energy_Bin_Pos_866 <= s_Energy_Bin_Pos_866;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_866 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_866;   
  
 Energy_Bin_Pos_867 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_867   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_867 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E867_C1_L_Pos and PEAK_C1_Pos <= s_E867_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_867 <= s_Energy_Bin_Pos_867 +'1';
		 Energy_Bin_Pos_Rdy_867 <= '1';
		else
		 s_Energy_Bin_Pos_867 <= s_Energy_Bin_Pos_867;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_867 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_867;   
  
  Energy_Bin_Pos_868 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_868   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_868 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E868_C1_L_Pos and PEAK_C1_Pos <= s_E868_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_868 <= s_Energy_Bin_Pos_868 +'1';
		 Energy_Bin_Pos_Rdy_868 <= '1';
		else
		 s_Energy_Bin_Pos_868 <= s_Energy_Bin_Pos_868;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_868 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_868;   
  
  Energy_Bin_Pos_869 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_869   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_869 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E869_C1_L_Pos and PEAK_C1_Pos <= s_E869_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_869 <= s_Energy_Bin_Pos_869 +'1';
		 Energy_Bin_Pos_Rdy_869 <= '1';
		else
		 s_Energy_Bin_Pos_869 <= s_Energy_Bin_Pos_869;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_869 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_869;         
  
     Energy_Bin_Pos_870 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_870   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_870 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E870_C1_L_Pos and PEAK_C1_Pos <= s_E870_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_870 <= s_Energy_Bin_Pos_870 +'1';
		 Energy_Bin_Pos_Rdy_870 <= '1';
		else
		 s_Energy_Bin_Pos_870 <= s_Energy_Bin_Pos_870;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_870 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_870;    
  
  Energy_Bin_Pos_871 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_871   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_871 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E871_C1_L_Pos and PEAK_C1_Pos <= s_E871_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_871 <= s_Energy_Bin_Pos_871 +'1';
		 Energy_Bin_Pos_Rdy_871 <= '1';
		else
		 s_Energy_Bin_Pos_871 <= s_Energy_Bin_Pos_871;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_871 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_871;   
  
  Energy_Bin_Pos_872 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_872   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_872 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E872_C1_L_Pos and PEAK_C1_Pos <= s_E872_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_872 <= s_Energy_Bin_Pos_872 +'1';
		 Energy_Bin_Pos_Rdy_872 <= '1';
		else
		 s_Energy_Bin_Pos_872 <= s_Energy_Bin_Pos_872;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_872 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_872;   
  
  Energy_Bin_Pos_873 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_873   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_873 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E873_C1_L_Pos and PEAK_C1_Pos <= s_E873_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_873 <= s_Energy_Bin_Pos_873 +'1';
		 Energy_Bin_Pos_Rdy_873 <= '1';
		else
		 s_Energy_Bin_Pos_873 <= s_Energy_Bin_Pos_873;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_873 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_873;   
  
  Energy_Bin_Pos_874 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_874   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_874 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E874_C1_L_Pos and PEAK_C1_Pos <= s_E874_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_874 <= s_Energy_Bin_Pos_874 +'1';
		 Energy_Bin_Pos_Rdy_874 <= '1';
		else
		 s_Energy_Bin_Pos_874 <= s_Energy_Bin_Pos_874;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_874 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_874;   
 
 
  Energy_Bin_Pos_875 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_875   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_875 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E875_C1_L_Pos and PEAK_C1_Pos <= s_E875_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_875 <= s_Energy_Bin_Pos_875 +'1';
		 Energy_Bin_Pos_Rdy_875 <= '1';
		else
		 s_Energy_Bin_Pos_875 <= s_Energy_Bin_Pos_875;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_875 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_875;  
 
  
  Energy_Bin_Pos_876 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_876   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_876 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E876_C1_L_Pos and PEAK_C1_Pos <= s_E876_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_876 <= s_Energy_Bin_Pos_876 +'1';
		 Energy_Bin_Pos_Rdy_876 <= '1';
		else
		 s_Energy_Bin_Pos_876 <= s_Energy_Bin_Pos_876;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_876 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_876;   
  
 Energy_Bin_Pos_877 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_877   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_877 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E877_C1_L_Pos and PEAK_C1_Pos <= s_E877_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_877 <= s_Energy_Bin_Pos_877 +'1';
		 Energy_Bin_Pos_Rdy_877 <= '1';
		else
		 s_Energy_Bin_Pos_877 <= s_Energy_Bin_Pos_877;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_877 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_877;   
  
  Energy_Bin_Pos_878 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_878   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_878 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E878_C1_L_Pos and PEAK_C1_Pos <= s_E878_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_878 <= s_Energy_Bin_Pos_878 +'1';
		 Energy_Bin_Pos_Rdy_878 <= '1';
		else
		 s_Energy_Bin_Pos_878 <= s_Energy_Bin_Pos_878;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_878 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_878;   
  
  Energy_Bin_Pos_879 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_879   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_879 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E879_C1_L_Pos and PEAK_C1_Pos <= s_E879_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_879 <= s_Energy_Bin_Pos_879 +'1';
		 Energy_Bin_Pos_Rdy_879 <= '1';
		else
		 s_Energy_Bin_Pos_879 <= s_Energy_Bin_Pos_879;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_879 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_879;       
  
     Energy_Bin_Pos_880 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_880   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_880 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E880_C1_L_Pos and PEAK_C1_Pos <= s_E880_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_880 <= s_Energy_Bin_Pos_880 +'1';
		 Energy_Bin_Pos_Rdy_880 <= '1';
		else
		 s_Energy_Bin_Pos_880 <= s_Energy_Bin_Pos_880;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_880 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_880;    
  
  Energy_Bin_Pos_881 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_881   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_881 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E881_C1_L_Pos and PEAK_C1_Pos <= s_E881_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_881 <= s_Energy_Bin_Pos_881 +'1';
		 Energy_Bin_Pos_Rdy_881 <= '1';
		else
		 s_Energy_Bin_Pos_881 <= s_Energy_Bin_Pos_881;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_881 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_881;   
  
  Energy_Bin_Pos_882 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_882   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_882 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E882_C1_L_Pos and PEAK_C1_Pos <= s_E882_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_882 <= s_Energy_Bin_Pos_882 +'1';
		 Energy_Bin_Pos_Rdy_882 <= '1';
		else
		 s_Energy_Bin_Pos_882 <= s_Energy_Bin_Pos_882;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_882 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_882;   
  
  Energy_Bin_Pos_883 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_883   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_883 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E883_C1_L_Pos and PEAK_C1_Pos <= s_E883_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_883 <= s_Energy_Bin_Pos_883 +'1';
		 Energy_Bin_Pos_Rdy_883 <= '1';
		else
		 s_Energy_Bin_Pos_883 <= s_Energy_Bin_Pos_883;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_883 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_883;   
  
  Energy_Bin_Pos_884 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_884   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_884 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E884_C1_L_Pos and PEAK_C1_Pos <= s_E884_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_884 <= s_Energy_Bin_Pos_884 +'1';
		 Energy_Bin_Pos_Rdy_884 <= '1';
		else
		 s_Energy_Bin_Pos_884 <= s_Energy_Bin_Pos_884;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_884 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_884;   
 
 
  Energy_Bin_Pos_885 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_885   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_885 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E885_C1_L_Pos and PEAK_C1_Pos <= s_E885_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_885 <= s_Energy_Bin_Pos_885 +'1';
		 Energy_Bin_Pos_Rdy_885 <= '1';
		else
		 s_Energy_Bin_Pos_885 <= s_Energy_Bin_Pos_885;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_885 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_885;  
 
  
  Energy_Bin_Pos_886 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_886   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_886 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E886_C1_L_Pos and PEAK_C1_Pos <= s_E886_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_886 <= s_Energy_Bin_Pos_886 +'1';
		 Energy_Bin_Pos_Rdy_886 <= '1';
		else
		 s_Energy_Bin_Pos_886 <= s_Energy_Bin_Pos_886;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_886 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_886;   
  
 Energy_Bin_Pos_887 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_887   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_887 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E887_C1_L_Pos and PEAK_C1_Pos <= s_E887_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_887 <= s_Energy_Bin_Pos_887 +'1';
		 Energy_Bin_Pos_Rdy_887 <= '1';
		else
		 s_Energy_Bin_Pos_887 <= s_Energy_Bin_Pos_887;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_887 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_887;   
  
  Energy_Bin_Pos_888 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_888   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_888 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E888_C1_L_Pos and PEAK_C1_Pos <= s_E888_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_888 <= s_Energy_Bin_Pos_888 +'1';
		 Energy_Bin_Pos_Rdy_888 <= '1';
		else
		 s_Energy_Bin_Pos_888 <= s_Energy_Bin_Pos_888;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_888 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_888;   
  
  Energy_Bin_Pos_889 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_889   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_889 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E889_C1_L_Pos and PEAK_C1_Pos <= s_E889_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_889 <= s_Energy_Bin_Pos_889 +'1';
		 Energy_Bin_Pos_Rdy_889 <= '1';
		else
		 s_Energy_Bin_Pos_889 <= s_Energy_Bin_Pos_889;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_889 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_889;      
  
     Energy_Bin_Pos_890 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_890   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_890 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E890_C1_L_Pos and PEAK_C1_Pos <= s_E890_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_890 <= s_Energy_Bin_Pos_890 +'1';
		 Energy_Bin_Pos_Rdy_890 <= '1';
		else
		 s_Energy_Bin_Pos_890 <= s_Energy_Bin_Pos_890;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_890 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_890;    
  
  Energy_Bin_Pos_891 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_891   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_891 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E891_C1_L_Pos and PEAK_C1_Pos <= s_E891_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_891 <= s_Energy_Bin_Pos_891 +'1';
		 Energy_Bin_Pos_Rdy_891 <= '1';
		else
		 s_Energy_Bin_Pos_891 <= s_Energy_Bin_Pos_891;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_891 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_891;   
  
  Energy_Bin_Pos_892 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_892   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_892 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E892_C1_L_Pos and PEAK_C1_Pos <= s_E892_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_892 <= s_Energy_Bin_Pos_892 +'1';
		 Energy_Bin_Pos_Rdy_892 <= '1';
		else
		 s_Energy_Bin_Pos_892 <= s_Energy_Bin_Pos_892;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_892 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_892;   
  
  Energy_Bin_Pos_893 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_893   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_893 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E893_C1_L_Pos and PEAK_C1_Pos <= s_E893_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_893 <= s_Energy_Bin_Pos_893 +'1';
		 Energy_Bin_Pos_Rdy_893 <= '1';
		else
		 s_Energy_Bin_Pos_893 <= s_Energy_Bin_Pos_893;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_893 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_893;   
  
  Energy_Bin_Pos_894 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_894   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_894 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E894_C1_L_Pos and PEAK_C1_Pos <= s_E894_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_894 <= s_Energy_Bin_Pos_894 +'1';
		 Energy_Bin_Pos_Rdy_894 <= '1';
		else
		 s_Energy_Bin_Pos_894 <= s_Energy_Bin_Pos_894;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_894 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_894;   
 
 
  Energy_Bin_Pos_895 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_895   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_895 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E895_C1_L_Pos and PEAK_C1_Pos <= s_E895_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_895 <= s_Energy_Bin_Pos_895 +'1';
		 Energy_Bin_Pos_Rdy_895 <= '1';
		else
		 s_Energy_Bin_Pos_895 <= s_Energy_Bin_Pos_895;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_895 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_895;  
 
  
  Energy_Bin_Pos_896 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_896   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_896 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E896_C1_L_Pos and PEAK_C1_Pos <= s_E896_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_896 <= s_Energy_Bin_Pos_896 +'1';
		 Energy_Bin_Pos_Rdy_896 <= '1';
		else
		 s_Energy_Bin_Pos_896 <= s_Energy_Bin_Pos_896;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_896 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_896;   
  
 Energy_Bin_Pos_897 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_897   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_897 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E897_C1_L_Pos and PEAK_C1_Pos <= s_E897_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_897 <= s_Energy_Bin_Pos_897 +'1';
		 Energy_Bin_Pos_Rdy_897 <= '1';
		else
		 s_Energy_Bin_Pos_897 <= s_Energy_Bin_Pos_897;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_897 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_897;   
  
  Energy_Bin_Pos_898 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_898   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_898 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E898_C1_L_Pos and PEAK_C1_Pos <= s_E898_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_898 <= s_Energy_Bin_Pos_898 +'1';
		 Energy_Bin_Pos_Rdy_898 <= '1';
		else
		 s_Energy_Bin_Pos_898 <= s_Energy_Bin_Pos_898;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_898 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_898;   
  
  Energy_Bin_Pos_899 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_899   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_899 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E899_C1_L_Pos and PEAK_C1_Pos <= s_E899_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_899 <= s_Energy_Bin_Pos_899 +'1';
		 Energy_Bin_Pos_Rdy_899 <= '1';
		else
		 s_Energy_Bin_Pos_899 <= s_Energy_Bin_Pos_899;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_899 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_899;   

    Energy_Bin_Pos_900 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_900   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_900 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E900_C1_L_Pos and PEAK_C1_Pos <= s_E900_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_900 <= s_Energy_Bin_Pos_900 +'1';
		 Energy_Bin_Pos_Rdy_900 <= '1';
		else
		 s_Energy_Bin_Pos_900 <= s_Energy_Bin_Pos_900;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_900 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_900;    
  
  Energy_Bin_Pos_901 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_901   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_901 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E901_C1_L_Pos and PEAK_C1_Pos <= s_E901_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_901 <= s_Energy_Bin_Pos_901 +'1';
		 Energy_Bin_Pos_Rdy_901 <= '1';
		else
		 s_Energy_Bin_Pos_901 <= s_Energy_Bin_Pos_901;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_901 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_901;   
  
  Energy_Bin_Pos_902 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_902   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_902 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E902_C1_L_Pos and PEAK_C1_Pos <= s_E902_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_902 <= s_Energy_Bin_Pos_902 +'1';
		 Energy_Bin_Pos_Rdy_902 <= '1';
		else
		 s_Energy_Bin_Pos_902 <= s_Energy_Bin_Pos_902;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_902 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_902;   
  
  Energy_Bin_Pos_903 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_903   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_903 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E903_C1_L_Pos and PEAK_C1_Pos <= s_E903_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_903 <= s_Energy_Bin_Pos_903 +'1';
		 Energy_Bin_Pos_Rdy_903 <= '1';
		else
		 s_Energy_Bin_Pos_903 <= s_Energy_Bin_Pos_903;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_903 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_903;   
  
  Energy_Bin_Pos_904 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_904   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_904 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E904_C1_L_Pos and PEAK_C1_Pos <= s_E904_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_904 <= s_Energy_Bin_Pos_904 +'1';
		 Energy_Bin_Pos_Rdy_904 <= '1';
		else
		 s_Energy_Bin_Pos_904 <= s_Energy_Bin_Pos_904;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_904 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_904;   
 
 
  Energy_Bin_Pos_905 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_905   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_905 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E905_C1_L_Pos and PEAK_C1_Pos <= s_E905_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_905 <= s_Energy_Bin_Pos_905 +'1';
		 Energy_Bin_Pos_Rdy_905 <= '1';
		else
		 s_Energy_Bin_Pos_905 <= s_Energy_Bin_Pos_905;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_905 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_905;  
 
  
  Energy_Bin_Pos_906 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_906   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_906 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E906_C1_L_Pos and PEAK_C1_Pos <= s_E906_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_906 <= s_Energy_Bin_Pos_906 +'1';
		 Energy_Bin_Pos_Rdy_906 <= '1';
		else
		 s_Energy_Bin_Pos_906 <= s_Energy_Bin_Pos_906;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_906 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_906;   
  
 Energy_Bin_Pos_907 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_907   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_907 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E907_C1_L_Pos and PEAK_C1_Pos <= s_E907_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_907 <= s_Energy_Bin_Pos_907 +'1';
		 Energy_Bin_Pos_Rdy_907 <= '1';
		else
		 s_Energy_Bin_Pos_907 <= s_Energy_Bin_Pos_907;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_907 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_907;   
  
  Energy_Bin_Pos_908 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_908   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_908 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E908_C1_L_Pos and PEAK_C1_Pos <= s_E908_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_908 <= s_Energy_Bin_Pos_908 +'1';
		 Energy_Bin_Pos_Rdy_908 <= '1';
		else
		 s_Energy_Bin_Pos_908 <= s_Energy_Bin_Pos_908;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_908 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_908;   
  
  Energy_Bin_Pos_909 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_909   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_909 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E909_C1_L_Pos and PEAK_C1_Pos <= s_E909_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_909 <= s_Energy_Bin_Pos_909 +'1';
		 Energy_Bin_Pos_Rdy_909 <= '1';
		else
		 s_Energy_Bin_Pos_909 <= s_Energy_Bin_Pos_909;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_909 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_909;      
  
     Energy_Bin_Pos_910 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_910   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_910 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E910_C1_L_Pos and PEAK_C1_Pos <= s_E910_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_910 <= s_Energy_Bin_Pos_910 +'1';
		 Energy_Bin_Pos_Rdy_910 <= '1';
		else
		 s_Energy_Bin_Pos_910 <= s_Energy_Bin_Pos_910;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_910 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_910;    
  
  Energy_Bin_Pos_911 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_911   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_911 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E911_C1_L_Pos and PEAK_C1_Pos <= s_E911_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_911 <= s_Energy_Bin_Pos_911 +'1';
		 Energy_Bin_Pos_Rdy_911 <= '1';
		else
		 s_Energy_Bin_Pos_911 <= s_Energy_Bin_Pos_911;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_911 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_911;   
  
  Energy_Bin_Pos_912 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_912   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_912 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E912_C1_L_Pos and PEAK_C1_Pos <= s_E912_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_912 <= s_Energy_Bin_Pos_912 +'1';
		 Energy_Bin_Pos_Rdy_912 <= '1';
		else
		 s_Energy_Bin_Pos_912 <= s_Energy_Bin_Pos_912;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_912 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_912;   
  
  Energy_Bin_Pos_913 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_913   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_913 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E913_C1_L_Pos and PEAK_C1_Pos <= s_E913_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_913 <= s_Energy_Bin_Pos_913 +'1';
		 Energy_Bin_Pos_Rdy_913 <= '1';
		else
		 s_Energy_Bin_Pos_913 <= s_Energy_Bin_Pos_913;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_913 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_913;   
  
  Energy_Bin_Pos_914 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_914   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_914 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E914_C1_L_Pos and PEAK_C1_Pos <= s_E914_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_914 <= s_Energy_Bin_Pos_914 +'1';
		 Energy_Bin_Pos_Rdy_914 <= '1';
		else
		 s_Energy_Bin_Pos_914 <= s_Energy_Bin_Pos_914;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_914 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_914;   
 
 
  Energy_Bin_Pos_915 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_915   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_915 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E915_C1_L_Pos and PEAK_C1_Pos <= s_E915_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_915 <= s_Energy_Bin_Pos_915 +'1';
		 Energy_Bin_Pos_Rdy_915 <= '1';
		else
		 s_Energy_Bin_Pos_915 <= s_Energy_Bin_Pos_915;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_915 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_915;  
 
  
  Energy_Bin_Pos_916 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_916   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_916 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E916_C1_L_Pos and PEAK_C1_Pos <= s_E916_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_916 <= s_Energy_Bin_Pos_916 +'1';
		 Energy_Bin_Pos_Rdy_916 <= '1';
		else
		 s_Energy_Bin_Pos_916 <= s_Energy_Bin_Pos_916;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_916 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_916;   
  
 Energy_Bin_Pos_917 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_917   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_917 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E917_C1_L_Pos and PEAK_C1_Pos <= s_E917_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_917 <= s_Energy_Bin_Pos_917 +'1';
		 Energy_Bin_Pos_Rdy_917 <= '1';
		else
		 s_Energy_Bin_Pos_917 <= s_Energy_Bin_Pos_917;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_917 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_917;   
  
  Energy_Bin_Pos_918 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_918   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_918 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E918_C1_L_Pos and PEAK_C1_Pos <= s_E918_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_918 <= s_Energy_Bin_Pos_918 +'1';
		 Energy_Bin_Pos_Rdy_918 <= '1';
		else
		 s_Energy_Bin_Pos_918 <= s_Energy_Bin_Pos_918;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_918 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_918;   
  
  Energy_Bin_Pos_919 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_919   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_919 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E919_C1_L_Pos and PEAK_C1_Pos <= s_E919_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_919 <= s_Energy_Bin_Pos_919 +'1';
		 Energy_Bin_Pos_Rdy_919 <= '1';
		else
		 s_Energy_Bin_Pos_919 <= s_Energy_Bin_Pos_919;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_919 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_919;       
  
     Energy_Bin_Pos_920 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_920   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_920 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E920_C1_L_Pos and PEAK_C1_Pos <= s_E920_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_920 <= s_Energy_Bin_Pos_920 +'1';
		 Energy_Bin_Pos_Rdy_920 <= '1';
		else
		 s_Energy_Bin_Pos_920 <= s_Energy_Bin_Pos_920;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_920 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_920;    
  
  Energy_Bin_Pos_921 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_921   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_921 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E921_C1_L_Pos and PEAK_C1_Pos <= s_E921_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_921 <= s_Energy_Bin_Pos_921 +'1';
		 Energy_Bin_Pos_Rdy_921 <= '1';
		else
		 s_Energy_Bin_Pos_921 <= s_Energy_Bin_Pos_921;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_921 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_921;   
  
  Energy_Bin_Pos_922 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_922   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_922 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E922_C1_L_Pos and PEAK_C1_Pos <= s_E922_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_922 <= s_Energy_Bin_Pos_922 +'1';
		 Energy_Bin_Pos_Rdy_922 <= '1';
		else
		 s_Energy_Bin_Pos_922 <= s_Energy_Bin_Pos_922;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_922 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_922;   
  
  Energy_Bin_Pos_923 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_923   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_923 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E923_C1_L_Pos and PEAK_C1_Pos <= s_E923_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_923 <= s_Energy_Bin_Pos_923 +'1';
		 Energy_Bin_Pos_Rdy_923 <= '1';
		else
		 s_Energy_Bin_Pos_923 <= s_Energy_Bin_Pos_923;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_923 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_923;   
  
  Energy_Bin_Pos_924 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_924   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_924 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E924_C1_L_Pos and PEAK_C1_Pos <= s_E924_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_924 <= s_Energy_Bin_Pos_924 +'1';
		 Energy_Bin_Pos_Rdy_924 <= '1';
		else
		 s_Energy_Bin_Pos_924 <= s_Energy_Bin_Pos_924;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_924 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_924;   
 
 
  Energy_Bin_Pos_925 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_925   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_925 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E925_C1_L_Pos and PEAK_C1_Pos <= s_E925_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_925 <= s_Energy_Bin_Pos_925 +'1';
		 Energy_Bin_Pos_Rdy_925 <= '1';
		else
		 s_Energy_Bin_Pos_925 <= s_Energy_Bin_Pos_925;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_925 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_925;  
 
  
  Energy_Bin_Pos_926 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_926   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_926 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E926_C1_L_Pos and PEAK_C1_Pos <= s_E926_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_926 <= s_Energy_Bin_Pos_926 +'1';
		 Energy_Bin_Pos_Rdy_926 <= '1';
		else
		 s_Energy_Bin_Pos_926 <= s_Energy_Bin_Pos_926;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_926 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_926;   
  
 Energy_Bin_Pos_927 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_927   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_927 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E927_C1_L_Pos and PEAK_C1_Pos <= s_E927_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_927 <= s_Energy_Bin_Pos_927 +'1';
		 Energy_Bin_Pos_Rdy_927 <= '1';
		else
		 s_Energy_Bin_Pos_927 <= s_Energy_Bin_Pos_927;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_927 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_927;   
  
  Energy_Bin_Pos_928 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_928   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_928 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E928_C1_L_Pos and PEAK_C1_Pos <= s_E928_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_928 <= s_Energy_Bin_Pos_928 +'1';
		 Energy_Bin_Pos_Rdy_928 <= '1';
		else
		 s_Energy_Bin_Pos_928 <= s_Energy_Bin_Pos_928;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_928 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_928;   
  
  Energy_Bin_Pos_929 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_929   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_929 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E929_C1_L_Pos and PEAK_C1_Pos <= s_E929_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_929 <= s_Energy_Bin_Pos_929 +'1';
		 Energy_Bin_Pos_Rdy_929 <= '1';
		else
		 s_Energy_Bin_Pos_929 <= s_Energy_Bin_Pos_929;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_929 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_929;        
  
     Energy_Bin_Pos_930 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_930   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_930 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E930_C1_L_Pos and PEAK_C1_Pos <= s_E930_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_930 <= s_Energy_Bin_Pos_930 +'1';
		 Energy_Bin_Pos_Rdy_930 <= '1';
		else
		 s_Energy_Bin_Pos_930 <= s_Energy_Bin_Pos_930;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_930 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_930;    
  
  Energy_Bin_Pos_931 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_931   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_931 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E931_C1_L_Pos and PEAK_C1_Pos <= s_E931_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_931 <= s_Energy_Bin_Pos_931 +'1';
		 Energy_Bin_Pos_Rdy_931 <= '1';
		else
		 s_Energy_Bin_Pos_931 <= s_Energy_Bin_Pos_931;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_931 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_931;   
  
  Energy_Bin_Pos_932 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_932   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_932 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E932_C1_L_Pos and PEAK_C1_Pos <= s_E932_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_932 <= s_Energy_Bin_Pos_932 +'1';
		 Energy_Bin_Pos_Rdy_932 <= '1';
		else
		 s_Energy_Bin_Pos_932 <= s_Energy_Bin_Pos_932;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_932 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_932;   
  
  Energy_Bin_Pos_933 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_933   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_933 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E933_C1_L_Pos and PEAK_C1_Pos <= s_E933_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_933 <= s_Energy_Bin_Pos_933 +'1';
		 Energy_Bin_Pos_Rdy_933 <= '1';
		else
		 s_Energy_Bin_Pos_933 <= s_Energy_Bin_Pos_933;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_933 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_933;   
  
  Energy_Bin_Pos_934 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_934   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_934 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E934_C1_L_Pos and PEAK_C1_Pos <= s_E934_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_934 <= s_Energy_Bin_Pos_934 +'1';
		 Energy_Bin_Pos_Rdy_934 <= '1';
		else
		 s_Energy_Bin_Pos_934 <= s_Energy_Bin_Pos_934;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_934 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_934;   
 
 
  Energy_Bin_Pos_935 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_935   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_935 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E935_C1_L_Pos and PEAK_C1_Pos <= s_E935_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_935 <= s_Energy_Bin_Pos_935 +'1';
		 Energy_Bin_Pos_Rdy_935 <= '1';
		else
		 s_Energy_Bin_Pos_935 <= s_Energy_Bin_Pos_935;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_935 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_935;  
 
  
  Energy_Bin_Pos_936 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_936   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_936 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E936_C1_L_Pos and PEAK_C1_Pos <= s_E936_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_936 <= s_Energy_Bin_Pos_936 +'1';
		 Energy_Bin_Pos_Rdy_936 <= '1';
		else
		 s_Energy_Bin_Pos_936 <= s_Energy_Bin_Pos_936;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_936 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_936;   
  
 Energy_Bin_Pos_937 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_937   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_937 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E937_C1_L_Pos and PEAK_C1_Pos <= s_E937_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_937 <= s_Energy_Bin_Pos_937 +'1';
		 Energy_Bin_Pos_Rdy_937 <= '1';
		else
		 s_Energy_Bin_Pos_937 <= s_Energy_Bin_Pos_937;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_937 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_937;   
  
  Energy_Bin_Pos_938 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_938   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_938 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E938_C1_L_Pos and PEAK_C1_Pos <= s_E938_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_938 <= s_Energy_Bin_Pos_938 +'1';
		 Energy_Bin_Pos_Rdy_938 <= '1';
		else
		 s_Energy_Bin_Pos_938 <= s_Energy_Bin_Pos_938;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_938 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_938;   
  
  Energy_Bin_Pos_939 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_939   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_939 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E939_C1_L_Pos and PEAK_C1_Pos <= s_E939_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_939 <= s_Energy_Bin_Pos_939 +'1';
		 Energy_Bin_Pos_Rdy_939 <= '1';
		else
		 s_Energy_Bin_Pos_939 <= s_Energy_Bin_Pos_939;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_939 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_939;         
  
     Energy_Bin_Pos_940 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_940   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_940 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E940_C1_L_Pos and PEAK_C1_Pos <= s_E940_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_940 <= s_Energy_Bin_Pos_940 +'1';
		 Energy_Bin_Pos_Rdy_940 <= '1';
		else
		 s_Energy_Bin_Pos_940 <= s_Energy_Bin_Pos_940;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_940 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_940;    
  
  Energy_Bin_Pos_941 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_941   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_941 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E941_C1_L_Pos and PEAK_C1_Pos <= s_E941_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_941 <= s_Energy_Bin_Pos_941 +'1';
		 Energy_Bin_Pos_Rdy_941 <= '1';
		else
		 s_Energy_Bin_Pos_941 <= s_Energy_Bin_Pos_941;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_941 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_941;   
  
  Energy_Bin_Pos_942 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_942   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_942 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E942_C1_L_Pos and PEAK_C1_Pos <= s_E942_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_942 <= s_Energy_Bin_Pos_942 +'1';
		 Energy_Bin_Pos_Rdy_942 <= '1';
		else
		 s_Energy_Bin_Pos_942 <= s_Energy_Bin_Pos_942;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_942 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_942;   
  
  Energy_Bin_Pos_943 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_943   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_943 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E943_C1_L_Pos and PEAK_C1_Pos <= s_E943_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_943 <= s_Energy_Bin_Pos_943 +'1';
		 Energy_Bin_Pos_Rdy_943 <= '1';
		else
		 s_Energy_Bin_Pos_943 <= s_Energy_Bin_Pos_943;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_943 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_943;   
  
  Energy_Bin_Pos_944 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_944   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_944 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E944_C1_L_Pos and PEAK_C1_Pos <= s_E944_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_944 <= s_Energy_Bin_Pos_944 +'1';
		 Energy_Bin_Pos_Rdy_944 <= '1';
		else
		 s_Energy_Bin_Pos_944 <= s_Energy_Bin_Pos_944;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_944 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_944;   
 
 
  Energy_Bin_Pos_945 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_945   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_945 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E945_C1_L_Pos and PEAK_C1_Pos <= s_E945_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_945 <= s_Energy_Bin_Pos_945 +'1';
		 Energy_Bin_Pos_Rdy_945 <= '1';
		else
		 s_Energy_Bin_Pos_945 <= s_Energy_Bin_Pos_945;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_945 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_945;  
 
  
  Energy_Bin_Pos_946 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_946   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_946 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E946_C1_L_Pos and PEAK_C1_Pos <= s_E946_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_946 <= s_Energy_Bin_Pos_946 +'1';
		 Energy_Bin_Pos_Rdy_946 <= '1';
		else
		 s_Energy_Bin_Pos_946 <= s_Energy_Bin_Pos_946;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_946 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_946;   
  
 Energy_Bin_Pos_947 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_947   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_947 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E947_C1_L_Pos and PEAK_C1_Pos <= s_E947_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_947 <= s_Energy_Bin_Pos_947 +'1';
		 Energy_Bin_Pos_Rdy_947 <= '1';
		else
		 s_Energy_Bin_Pos_947 <= s_Energy_Bin_Pos_947;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_947 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_947;   
  
  Energy_Bin_Pos_948 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_948   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_948 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E948_C1_L_Pos and PEAK_C1_Pos <= s_E948_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_948 <= s_Energy_Bin_Pos_948 +'1';
		 Energy_Bin_Pos_Rdy_948 <= '1';
		else
		 s_Energy_Bin_Pos_948 <= s_Energy_Bin_Pos_948;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_948 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_948;   
  
  Energy_Bin_Pos_949 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_949   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_949 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E949_C1_L_Pos and PEAK_C1_Pos <= s_E949_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_949 <= s_Energy_Bin_Pos_949 +'1';
		 Energy_Bin_Pos_Rdy_949 <= '1';
		else
		 s_Energy_Bin_Pos_949 <= s_Energy_Bin_Pos_949;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_949 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_949;          
  
  
     Energy_Bin_Pos_950 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_950   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_950 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E950_C1_L_Pos and PEAK_C1_Pos <= s_E950_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_950 <= s_Energy_Bin_Pos_950 +'1';
		 Energy_Bin_Pos_Rdy_950 <= '1';
		else
		 s_Energy_Bin_Pos_950 <= s_Energy_Bin_Pos_950;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_950 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_950;    
  
  Energy_Bin_Pos_951 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_951   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_951 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E951_C1_L_Pos and PEAK_C1_Pos <= s_E951_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_951 <= s_Energy_Bin_Pos_951 +'1';
		 Energy_Bin_Pos_Rdy_951 <= '1';
		else
		 s_Energy_Bin_Pos_951 <= s_Energy_Bin_Pos_951;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_951 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_951;   
  
  Energy_Bin_Pos_952 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_952   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_952 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E952_C1_L_Pos and PEAK_C1_Pos <= s_E952_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_952 <= s_Energy_Bin_Pos_952 +'1';
		 Energy_Bin_Pos_Rdy_952 <= '1';
		else
		 s_Energy_Bin_Pos_952 <= s_Energy_Bin_Pos_952;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_952 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_952;   
  
  Energy_Bin_Pos_953 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_953   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_953 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E953_C1_L_Pos and PEAK_C1_Pos <= s_E953_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_953 <= s_Energy_Bin_Pos_953 +'1';
		 Energy_Bin_Pos_Rdy_953 <= '1';
		else
		 s_Energy_Bin_Pos_953 <= s_Energy_Bin_Pos_953;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_953 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_953;   
  
  Energy_Bin_Pos_954 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_954   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_954 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E954_C1_L_Pos and PEAK_C1_Pos <= s_E954_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_954 <= s_Energy_Bin_Pos_954 +'1';
		 Energy_Bin_Pos_Rdy_954 <= '1';
		else
		 s_Energy_Bin_Pos_954 <= s_Energy_Bin_Pos_954;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_954 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_954;   
 
 
  Energy_Bin_Pos_955 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_955   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_955 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E955_C1_L_Pos and PEAK_C1_Pos <= s_E955_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_955 <= s_Energy_Bin_Pos_955 +'1';
		 Energy_Bin_Pos_Rdy_955 <= '1';
		else
		 s_Energy_Bin_Pos_955 <= s_Energy_Bin_Pos_955;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_955 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_955;  
 
  
  Energy_Bin_Pos_956 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_956   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_956 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E956_C1_L_Pos and PEAK_C1_Pos <= s_E956_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_956 <= s_Energy_Bin_Pos_956 +'1';
		 Energy_Bin_Pos_Rdy_956 <= '1';
		else
		 s_Energy_Bin_Pos_956 <= s_Energy_Bin_Pos_956;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_956 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_956;   
  
 Energy_Bin_Pos_957 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_957   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_957 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E957_C1_L_Pos and PEAK_C1_Pos <= s_E957_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_957 <= s_Energy_Bin_Pos_957 +'1';
		 Energy_Bin_Pos_Rdy_957 <= '1';
		else
		 s_Energy_Bin_Pos_957 <= s_Energy_Bin_Pos_957;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_957 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_957;   
  
  Energy_Bin_Pos_958 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_958   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_958 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E958_C1_L_Pos and PEAK_C1_Pos <= s_E958_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_958 <= s_Energy_Bin_Pos_958 +'1';
		 Energy_Bin_Pos_Rdy_958 <= '1';
		else
		 s_Energy_Bin_Pos_958 <= s_Energy_Bin_Pos_958;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_958 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_958;   
  
  Energy_Bin_Pos_959 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_959   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_959 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E959_C1_L_Pos and PEAK_C1_Pos <= s_E959_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_959 <= s_Energy_Bin_Pos_959 +'1';
		 Energy_Bin_Pos_Rdy_959 <= '1';
		else
		 s_Energy_Bin_Pos_959 <= s_Energy_Bin_Pos_959;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_959 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_959;           
  
     Energy_Bin_Pos_960 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_960   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_960 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E960_C1_L_Pos and PEAK_C1_Pos <= s_E960_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_960 <= s_Energy_Bin_Pos_960 +'1';
		 Energy_Bin_Pos_Rdy_960 <= '1';
		else
		 s_Energy_Bin_Pos_960 <= s_Energy_Bin_Pos_960;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_960 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_960;    
  
  Energy_Bin_Pos_961 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_961   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_961 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E961_C1_L_Pos and PEAK_C1_Pos <= s_E961_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_961 <= s_Energy_Bin_Pos_961 +'1';
		 Energy_Bin_Pos_Rdy_961 <= '1';
		else
		 s_Energy_Bin_Pos_961 <= s_Energy_Bin_Pos_961;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_961 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_961;   
  
  Energy_Bin_Pos_962 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_962   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_962 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E962_C1_L_Pos and PEAK_C1_Pos <= s_E962_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_962 <= s_Energy_Bin_Pos_962 +'1';
		 Energy_Bin_Pos_Rdy_962 <= '1';
		else
		 s_Energy_Bin_Pos_962 <= s_Energy_Bin_Pos_962;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_962 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_962;   
  
  Energy_Bin_Pos_963 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_963   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_963 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E963_C1_L_Pos and PEAK_C1_Pos <= s_E963_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_963 <= s_Energy_Bin_Pos_963 +'1';
		 Energy_Bin_Pos_Rdy_963 <= '1';
		else
		 s_Energy_Bin_Pos_963 <= s_Energy_Bin_Pos_963;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_963 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_963;   
  
  Energy_Bin_Pos_964 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_964   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_964 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E964_C1_L_Pos and PEAK_C1_Pos <= s_E964_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_964 <= s_Energy_Bin_Pos_964 +'1';
		 Energy_Bin_Pos_Rdy_964 <= '1';
		else
		 s_Energy_Bin_Pos_964 <= s_Energy_Bin_Pos_964;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_964 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_964;   
 
 
  Energy_Bin_Pos_965 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_965   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_965 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E965_C1_L_Pos and PEAK_C1_Pos <= s_E965_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_965 <= s_Energy_Bin_Pos_965 +'1';
		 Energy_Bin_Pos_Rdy_965 <= '1';
		else
		 s_Energy_Bin_Pos_965 <= s_Energy_Bin_Pos_965;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_965 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_965;  
 
  
  Energy_Bin_Pos_966 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_966   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_966 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E966_C1_L_Pos and PEAK_C1_Pos <= s_E966_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_966 <= s_Energy_Bin_Pos_966 +'1';
		 Energy_Bin_Pos_Rdy_966 <= '1';
		else
		 s_Energy_Bin_Pos_966 <= s_Energy_Bin_Pos_966;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_966 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_966;   
  
 Energy_Bin_Pos_967 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_967   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_967 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E967_C1_L_Pos and PEAK_C1_Pos <= s_E967_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_967 <= s_Energy_Bin_Pos_967 +'1';
		 Energy_Bin_Pos_Rdy_967 <= '1';
		else
		 s_Energy_Bin_Pos_967 <= s_Energy_Bin_Pos_967;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_967 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_967;   
  
  Energy_Bin_Pos_968 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_968   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_968 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E968_C1_L_Pos and PEAK_C1_Pos <= s_E968_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_968 <= s_Energy_Bin_Pos_968 +'1';
		 Energy_Bin_Pos_Rdy_968 <= '1';
		else
		 s_Energy_Bin_Pos_968 <= s_Energy_Bin_Pos_968;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_968 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_968;   
  
  Energy_Bin_Pos_969 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_969   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_969 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E969_C1_L_Pos and PEAK_C1_Pos <= s_E969_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_969 <= s_Energy_Bin_Pos_969 +'1';
		 Energy_Bin_Pos_Rdy_969 <= '1';
		else
		 s_Energy_Bin_Pos_969 <= s_Energy_Bin_Pos_969;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_969 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_969;         
  
     Energy_Bin_Pos_970 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_970   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_970 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E970_C1_L_Pos and PEAK_C1_Pos <= s_E970_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_970 <= s_Energy_Bin_Pos_970 +'1';
		 Energy_Bin_Pos_Rdy_970 <= '1';
		else
		 s_Energy_Bin_Pos_970 <= s_Energy_Bin_Pos_970;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_970 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_970;    
  
  Energy_Bin_Pos_971 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_971   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_971 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E971_C1_L_Pos and PEAK_C1_Pos <= s_E971_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_971 <= s_Energy_Bin_Pos_971 +'1';
		 Energy_Bin_Pos_Rdy_971 <= '1';
		else
		 s_Energy_Bin_Pos_971 <= s_Energy_Bin_Pos_971;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_971 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_971;   
  
  Energy_Bin_Pos_972 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_972   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_972 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E972_C1_L_Pos and PEAK_C1_Pos <= s_E972_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_972 <= s_Energy_Bin_Pos_972 +'1';
		 Energy_Bin_Pos_Rdy_972 <= '1';
		else
		 s_Energy_Bin_Pos_972 <= s_Energy_Bin_Pos_972;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_972 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_972;   
  
  Energy_Bin_Pos_973 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_973   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_973 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E973_C1_L_Pos and PEAK_C1_Pos <= s_E973_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_973 <= s_Energy_Bin_Pos_973 +'1';
		 Energy_Bin_Pos_Rdy_973 <= '1';
		else
		 s_Energy_Bin_Pos_973 <= s_Energy_Bin_Pos_973;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_973 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_973;   
  
  Energy_Bin_Pos_974 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_974   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_974 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E974_C1_L_Pos and PEAK_C1_Pos <= s_E974_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_974 <= s_Energy_Bin_Pos_974 +'1';
		 Energy_Bin_Pos_Rdy_974 <= '1';
		else
		 s_Energy_Bin_Pos_974 <= s_Energy_Bin_Pos_974;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_974 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_974;   
 
 
  Energy_Bin_Pos_975 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_975   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_975 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E975_C1_L_Pos and PEAK_C1_Pos <= s_E975_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_975 <= s_Energy_Bin_Pos_975 +'1';
		 Energy_Bin_Pos_Rdy_975 <= '1';
		else
		 s_Energy_Bin_Pos_975 <= s_Energy_Bin_Pos_975;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_975 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_975;  
 
  
  Energy_Bin_Pos_976 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_976   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_976 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E976_C1_L_Pos and PEAK_C1_Pos <= s_E976_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_976 <= s_Energy_Bin_Pos_976 +'1';
		 Energy_Bin_Pos_Rdy_976 <= '1';
		else
		 s_Energy_Bin_Pos_976 <= s_Energy_Bin_Pos_976;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_976 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_976;   
  
 Energy_Bin_Pos_977 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_977   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_977 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E977_C1_L_Pos and PEAK_C1_Pos <= s_E977_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_977 <= s_Energy_Bin_Pos_977 +'1';
		 Energy_Bin_Pos_Rdy_977 <= '1';
		else
		 s_Energy_Bin_Pos_977 <= s_Energy_Bin_Pos_977;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_977 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_977;   
  
  Energy_Bin_Pos_978 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_978   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_978 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E978_C1_L_Pos and PEAK_C1_Pos <= s_E978_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_978 <= s_Energy_Bin_Pos_978 +'1';
		 Energy_Bin_Pos_Rdy_978 <= '1';
		else
		 s_Energy_Bin_Pos_978 <= s_Energy_Bin_Pos_978;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_978 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_978;   
  
  Energy_Bin_Pos_979 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_979   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_979 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E979_C1_L_Pos and PEAK_C1_Pos <= s_E979_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_979 <= s_Energy_Bin_Pos_979 +'1';
		 Energy_Bin_Pos_Rdy_979 <= '1';
		else
		 s_Energy_Bin_Pos_979 <= s_Energy_Bin_Pos_979;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_979 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_979;       
  
     Energy_Bin_Pos_980 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_980   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_980 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E980_C1_L_Pos and PEAK_C1_Pos <= s_E980_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_980 <= s_Energy_Bin_Pos_980 +'1';
		 Energy_Bin_Pos_Rdy_980 <= '1';
		else
		 s_Energy_Bin_Pos_980 <= s_Energy_Bin_Pos_980;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_980 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_980;    
  
  Energy_Bin_Pos_981 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_981   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_981 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E981_C1_L_Pos and PEAK_C1_Pos <= s_E981_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_981 <= s_Energy_Bin_Pos_981 +'1';
		 Energy_Bin_Pos_Rdy_981 <= '1';
		else
		 s_Energy_Bin_Pos_981 <= s_Energy_Bin_Pos_981;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_981 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_981;   
  
  Energy_Bin_Pos_982 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_982   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_982 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E982_C1_L_Pos and PEAK_C1_Pos <= s_E982_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_982 <= s_Energy_Bin_Pos_982 +'1';
		 Energy_Bin_Pos_Rdy_982 <= '1';
		else
		 s_Energy_Bin_Pos_982 <= s_Energy_Bin_Pos_982;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_982 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_982;   
  
  Energy_Bin_Pos_983 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_983   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_983 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E983_C1_L_Pos and PEAK_C1_Pos <= s_E983_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_983 <= s_Energy_Bin_Pos_983 +'1';
		 Energy_Bin_Pos_Rdy_983 <= '1';
		else
		 s_Energy_Bin_Pos_983 <= s_Energy_Bin_Pos_983;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_983 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_983;   
  
  Energy_Bin_Pos_984 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_984   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_984 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E984_C1_L_Pos and PEAK_C1_Pos <= s_E984_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_984 <= s_Energy_Bin_Pos_984 +'1';
		 Energy_Bin_Pos_Rdy_984 <= '1';
		else
		 s_Energy_Bin_Pos_984 <= s_Energy_Bin_Pos_984;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_984 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_984;   
 
 
  Energy_Bin_Pos_985 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_985   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_985 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E985_C1_L_Pos and PEAK_C1_Pos <= s_E985_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_985 <= s_Energy_Bin_Pos_985 +'1';
		 Energy_Bin_Pos_Rdy_985 <= '1';
		else
		 s_Energy_Bin_Pos_985 <= s_Energy_Bin_Pos_985;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_985 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_985;  
 
  
  Energy_Bin_Pos_986 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_986   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_986 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E986_C1_L_Pos and PEAK_C1_Pos <= s_E986_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_986 <= s_Energy_Bin_Pos_986 +'1';
		 Energy_Bin_Pos_Rdy_986 <= '1';
		else
		 s_Energy_Bin_Pos_986 <= s_Energy_Bin_Pos_986;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_986 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_986;   
  
 Energy_Bin_Pos_987 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_987   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_987 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E987_C1_L_Pos and PEAK_C1_Pos <= s_E987_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_987 <= s_Energy_Bin_Pos_987 +'1';
		 Energy_Bin_Pos_Rdy_987 <= '1';
		else
		 s_Energy_Bin_Pos_987 <= s_Energy_Bin_Pos_987;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_987 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_987;   
  
  Energy_Bin_Pos_988 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_988   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_988 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E988_C1_L_Pos and PEAK_C1_Pos <= s_E988_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_988 <= s_Energy_Bin_Pos_988 +'1';
		 Energy_Bin_Pos_Rdy_988 <= '1';
		else
		 s_Energy_Bin_Pos_988 <= s_Energy_Bin_Pos_988;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_988 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_988;   
  
  Energy_Bin_Pos_989 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_989   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_989 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E989_C1_L_Pos and PEAK_C1_Pos <= s_E989_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_989 <= s_Energy_Bin_Pos_989 +'1';
		 Energy_Bin_Pos_Rdy_989 <= '1';
		else
		 s_Energy_Bin_Pos_989 <= s_Energy_Bin_Pos_989;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_989 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_989;      
  
     Energy_Bin_Pos_990 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_990   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_990 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E990_C1_L_Pos and PEAK_C1_Pos <= s_E990_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_990 <= s_Energy_Bin_Pos_990 +'1';
		 Energy_Bin_Pos_Rdy_990 <= '1';
		else
		 s_Energy_Bin_Pos_990 <= s_Energy_Bin_Pos_990;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_990 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_990;    
  
  Energy_Bin_Pos_991 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_991   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_991 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E991_C1_L_Pos and PEAK_C1_Pos <= s_E991_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_991 <= s_Energy_Bin_Pos_991 +'1';
		 Energy_Bin_Pos_Rdy_991 <= '1';
		else
		 s_Energy_Bin_Pos_991 <= s_Energy_Bin_Pos_991;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_991 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_991;   
  
  Energy_Bin_Pos_992 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_992   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_992 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E992_C1_L_Pos and PEAK_C1_Pos <= s_E992_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_992 <= s_Energy_Bin_Pos_992 +'1';
		 Energy_Bin_Pos_Rdy_992 <= '1';
		else
		 s_Energy_Bin_Pos_992 <= s_Energy_Bin_Pos_992;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_992 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_992;   
  
  Energy_Bin_Pos_993 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_993   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_993 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E993_C1_L_Pos and PEAK_C1_Pos <= s_E993_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_993 <= s_Energy_Bin_Pos_993 +'1';
		 Energy_Bin_Pos_Rdy_993 <= '1';
		else
		 s_Energy_Bin_Pos_993 <= s_Energy_Bin_Pos_993;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_993 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_993;   
  
  Energy_Bin_Pos_994 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_994   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_994 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E994_C1_L_Pos and PEAK_C1_Pos <= s_E994_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_994 <= s_Energy_Bin_Pos_994 +'1';
		 Energy_Bin_Pos_Rdy_994 <= '1';
		else
		 s_Energy_Bin_Pos_994 <= s_Energy_Bin_Pos_994;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_994 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_994;   
 
 
  Energy_Bin_Pos_995 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_995   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_995 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E995_C1_L_Pos and PEAK_C1_Pos <= s_E995_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_995 <= s_Energy_Bin_Pos_995 +'1';
		 Energy_Bin_Pos_Rdy_995 <= '1';
		else
		 s_Energy_Bin_Pos_995 <= s_Energy_Bin_Pos_995;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_995 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_995;  
 
  
  Energy_Bin_Pos_996 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_996   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_996 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E996_C1_L_Pos and PEAK_C1_Pos <= s_E996_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_996 <= s_Energy_Bin_Pos_996 +'1';
		 Energy_Bin_Pos_Rdy_996 <= '1';
		else
		 s_Energy_Bin_Pos_996 <= s_Energy_Bin_Pos_996;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_996 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_996;   
  
 Energy_Bin_Pos_997 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_997   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_997 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E997_C1_L_Pos and PEAK_C1_Pos <= s_E997_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_997 <= s_Energy_Bin_Pos_997 +'1';
		 Energy_Bin_Pos_Rdy_997 <= '1';
		else
		 s_Energy_Bin_Pos_997 <= s_Energy_Bin_Pos_997;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_997 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_997;   
  
  Energy_Bin_Pos_998 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_998   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_998 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E998_C1_L_Pos and PEAK_C1_Pos <= s_E998_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_998 <= s_Energy_Bin_Pos_998 +'1';
		 Energy_Bin_Pos_Rdy_998 <= '1';
		else
		 s_Energy_Bin_Pos_998 <= s_Energy_Bin_Pos_998;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_998 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_998;   
  
  Energy_Bin_Pos_999 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_999   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_999 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E999_C1_L_Pos and PEAK_C1_Pos <= s_E999_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_999 <= s_Energy_Bin_Pos_999 +'1';
		 Energy_Bin_Pos_Rdy_999 <= '1';
		else
		 s_Energy_Bin_Pos_999 <= s_Energy_Bin_Pos_999;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_999 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_999;   

    Energy_Bin_Pos_1000 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1000   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1000 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E1000_C1_L_Pos and PEAK_C1_Pos <= s_E1000_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1000 <= s_Energy_Bin_Pos_1000 +'1';
		 Energy_Bin_Pos_Rdy_1000 <= '1';
		else
		 s_Energy_Bin_Pos_1000 <= s_Energy_Bin_Pos_1000;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1000 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1000;    
  
  Energy_Bin_Pos_1001 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1001   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1001 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E1001_C1_L_Pos and PEAK_C1_Pos <= s_E1001_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1001 <= s_Energy_Bin_Pos_1001 +'1';
		 Energy_Bin_Pos_Rdy_1001 <= '1';
		else
		 s_Energy_Bin_Pos_1001 <= s_Energy_Bin_Pos_1001;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1001 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1001;   
  
  Energy_Bin_Pos_1002 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1002   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_1002 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E1002_C1_L_Pos and PEAK_C1_Pos <= s_E1002_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1002 <= s_Energy_Bin_Pos_1002 +'1';
		 Energy_Bin_Pos_Rdy_1002 <= '1';
		else
		 s_Energy_Bin_Pos_1002 <= s_Energy_Bin_Pos_1002;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1002 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1002;   
  
  Energy_Bin_Pos_1003 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1003   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_1003 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E1003_C1_L_Pos and PEAK_C1_Pos <= s_E1003_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1003 <= s_Energy_Bin_Pos_1003 +'1';
		 Energy_Bin_Pos_Rdy_1003 <= '1';
		else
		 s_Energy_Bin_Pos_1003 <= s_Energy_Bin_Pos_1003;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1003 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1003;   
  
  Energy_Bin_Pos_1004 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1004   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1004 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E1004_C1_L_Pos and PEAK_C1_Pos <= s_E1004_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1004 <= s_Energy_Bin_Pos_1004 +'1';
		 Energy_Bin_Pos_Rdy_1004 <= '1';
		else
		 s_Energy_Bin_Pos_1004 <= s_Energy_Bin_Pos_1004;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1004 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_1004;   
 
 
  Energy_Bin_Pos_1005 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1005   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1005 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E1005_C1_L_Pos and PEAK_C1_Pos <= s_E1005_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1005 <= s_Energy_Bin_Pos_1005 +'1';
		 Energy_Bin_Pos_Rdy_1005 <= '1';
		else
		 s_Energy_Bin_Pos_1005 <= s_Energy_Bin_Pos_1005;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1005 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_1005;  
 
  
  Energy_Bin_Pos_1006 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1006   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1006 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E1006_C1_L_Pos and PEAK_C1_Pos <= s_E1006_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1006 <= s_Energy_Bin_Pos_1006 +'1';
		 Energy_Bin_Pos_Rdy_1006 <= '1';
		else
		 s_Energy_Bin_Pos_1006 <= s_Energy_Bin_Pos_1006;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1006 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1006;   
  
 Energy_Bin_Pos_1007 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1007   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1007 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E1007_C1_L_Pos and PEAK_C1_Pos <= s_E1007_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1007 <= s_Energy_Bin_Pos_1007 +'1';
		 Energy_Bin_Pos_Rdy_1007 <= '1';
		else
		 s_Energy_Bin_Pos_1007 <= s_Energy_Bin_Pos_1007;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1007 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1007;   
  
  Energy_Bin_Pos_1008 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1008   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1008 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E1008_C1_L_Pos and PEAK_C1_Pos <= s_E1008_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1008 <= s_Energy_Bin_Pos_1008 +'1';
		 Energy_Bin_Pos_Rdy_1008 <= '1';
		else
		 s_Energy_Bin_Pos_1008 <= s_Energy_Bin_Pos_1008;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1008 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1008;   
  
  Energy_Bin_Pos_1009 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1009   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1009 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E1009_C1_L_Pos and PEAK_C1_Pos <= s_E1009_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1009 <= s_Energy_Bin_Pos_1009 +'1';
		 Energy_Bin_Pos_Rdy_1009 <= '1';
		else
		 s_Energy_Bin_Pos_1009 <= s_Energy_Bin_Pos_1009;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1009 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1009;      
  
     Energy_Bin_Pos_1010 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1010   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1010 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E1010_C1_L_Pos and PEAK_C1_Pos <= s_E1010_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1010 <= s_Energy_Bin_Pos_1010 +'1';
		 Energy_Bin_Pos_Rdy_1010 <= '1';
		else
		 s_Energy_Bin_Pos_1010 <= s_Energy_Bin_Pos_1010;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1010 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1010;    
  
  Energy_Bin_Pos_1011 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1011   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1011 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E1011_C1_L_Pos and PEAK_C1_Pos <= s_E1011_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1011 <= s_Energy_Bin_Pos_1011 +'1';
		 Energy_Bin_Pos_Rdy_1011 <= '1';
		else
		 s_Energy_Bin_Pos_1011 <= s_Energy_Bin_Pos_1011;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1011 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1011;   
  
  Energy_Bin_Pos_1012 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1012   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_1012 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E1012_C1_L_Pos and PEAK_C1_Pos <= s_E1012_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1012 <= s_Energy_Bin_Pos_1012 +'1';
		 Energy_Bin_Pos_Rdy_1012 <= '1';
		else
		 s_Energy_Bin_Pos_1012 <= s_Energy_Bin_Pos_1012;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1012 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1012;   
  
  Energy_Bin_Pos_1013 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1013   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_1013 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E1013_C1_L_Pos and PEAK_C1_Pos <= s_E1013_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1013 <= s_Energy_Bin_Pos_1013 +'1';
		 Energy_Bin_Pos_Rdy_1013 <= '1';
		else
		 s_Energy_Bin_Pos_1013 <= s_Energy_Bin_Pos_1013;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1013 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1013;   
  
  Energy_Bin_Pos_1014 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1014   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1014 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E1014_C1_L_Pos and PEAK_C1_Pos <= s_E1014_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1014 <= s_Energy_Bin_Pos_1014 +'1';
		 Energy_Bin_Pos_Rdy_1014 <= '1';
		else
		 s_Energy_Bin_Pos_1014 <= s_Energy_Bin_Pos_1014;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1014 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_1014;   
 
 
  Energy_Bin_Pos_1015 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1015   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1015 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E1015_C1_L_Pos and PEAK_C1_Pos <= s_E1015_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1015 <= s_Energy_Bin_Pos_1015 +'1';
		 Energy_Bin_Pos_Rdy_1015 <= '1';
		else
		 s_Energy_Bin_Pos_1015 <= s_Energy_Bin_Pos_1015;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1015 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_1015;  
 
  
  Energy_Bin_Pos_1016 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1016   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1016 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E1016_C1_L_Pos and PEAK_C1_Pos <= s_E1016_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1016 <= s_Energy_Bin_Pos_1016 +'1';
		 Energy_Bin_Pos_Rdy_1016 <= '1';
		else
		 s_Energy_Bin_Pos_1016 <= s_Energy_Bin_Pos_1016;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1016 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1016;   
  
 Energy_Bin_Pos_1017 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1017   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1017 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E1017_C1_L_Pos and PEAK_C1_Pos <= s_E1017_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1017 <= s_Energy_Bin_Pos_1017 +'1';
		 Energy_Bin_Pos_Rdy_1017 <= '1';
		else
		 s_Energy_Bin_Pos_1017 <= s_Energy_Bin_Pos_1017;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1017 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1017;   
  
  Energy_Bin_Pos_1018 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1018   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1018 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E1018_C1_L_Pos and PEAK_C1_Pos <= s_E1018_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1018 <= s_Energy_Bin_Pos_1018 +'1';
		 Energy_Bin_Pos_Rdy_1018 <= '1';
		else
		 s_Energy_Bin_Pos_1018 <= s_Energy_Bin_Pos_1018;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1018 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1018;   
  
  Energy_Bin_Pos_1019 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1019   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1019 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E1019_C1_L_Pos and PEAK_C1_Pos <= s_E1019_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1019 <= s_Energy_Bin_Pos_1019 +'1';
		 Energy_Bin_Pos_Rdy_1019 <= '1';
		else
		 s_Energy_Bin_Pos_1019 <= s_Energy_Bin_Pos_1019;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1019 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1019;       
  
     Energy_Bin_Pos_1020 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1020   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1020 <= '0';
      elsif(PEAK_FL_Ris_pos = '1' ) then
	  
	    if(PEAK_C1_Pos > s_E1020_C1_L_Pos and PEAK_C1_Pos <= s_E1020_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1020 <= s_Energy_Bin_Pos_1020 +'1';
		 Energy_Bin_Pos_Rdy_1020 <= '1';
		else
		 s_Energy_Bin_Pos_1020 <= s_Energy_Bin_Pos_1020;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1020 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1020;    
  
  Energy_Bin_Pos_1021 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1021   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1021 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E1021_C1_L_Pos and PEAK_C1_Pos <= s_E1021_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1021 <= s_Energy_Bin_Pos_1021 +'1';
		 Energy_Bin_Pos_Rdy_1021 <= '1';
		else
		 s_Energy_Bin_Pos_1021 <= s_Energy_Bin_Pos_1021;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1021 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1021;   
  
  Energy_Bin_Pos_1022 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1022   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_1022 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E1022_C1_L_Pos and PEAK_C1_Pos <= s_E1022_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1022 <= s_Energy_Bin_Pos_1022 +'1';
		 Energy_Bin_Pos_Rdy_1022 <= '1';
		else
		 s_Energy_Bin_Pos_1022 <= s_Energy_Bin_Pos_1022;
		end if;
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1022 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1022;   
  
  Energy_Bin_Pos_1023 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1023   <=  (others =>'0');
	    Energy_Bin_Pos_Rdy_1023 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E1023_C1_L_Pos and PEAK_C1_Pos <= s_E1023_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1023 <= s_Energy_Bin_Pos_1023 +'1';
		 Energy_Bin_Pos_Rdy_1023 <= '1';
		else
		 s_Energy_Bin_Pos_1023 <= s_Energy_Bin_Pos_1023;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1023 <= '0';
      end if;
    end if;
  end process  Energy_Bin_Pos_1023;   
  
  Energy_Bin_Pos_1024 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_1024   <=  (others =>'0');
		Energy_Bin_Pos_Rdy_1024 <= '0';
      elsif(PEAK_FL_Ris_pos = '1') then
	  
	    if(PEAK_C1_Pos > s_E1024_C1_L_Pos and PEAK_C1_Pos <= s_E1024_C1_H_Pos and Bin_OR_Pos = '0') then
         s_Energy_Bin_Pos_1024 <= s_Energy_Bin_Pos_1024 +'1';
		 Energy_Bin_Pos_Rdy_1024 <= '1';
		else
		 s_Energy_Bin_Pos_1024 <= s_Energy_Bin_Pos_1024;
		end if;
		
	  elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_1024 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_Pos_1024;   


  Energy_Bin_Pos_reject : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_Pos_reject   <=  (others =>'0');
        Energy_Bin_Pos_Rdy_reject <= '0';
      elsif(PEAK_FL_Ris_pos_s = '1' ) then
	    if(Energy_Bin_Pos_Rdy = '0') then
         s_Energy_Bin_Pos_reject <= s_Energy_Bin_Pos_reject +'1';
         Energy_Bin_Pos_Rdy_reject <= '1';
		else
		 s_Energy_Bin_Pos_reject <= s_Energy_Bin_Pos_reject;
		end if;
		
      elsif(Energy_Ris_Dis_Pos = '1') then
	    Energy_Bin_Pos_Rdy_reject <= '0';
      end if;
    end if;
 end process  Energy_Bin_Pos_reject;  
  
-- channel_1 negative energy bin
 Energy_Bin_1 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1   <=  (others =>'0');
		Energy_Bin_Rdy_1 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E1_C1_L and PEAK_C1 <= s_E1_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1 <= s_Energy_Bin_1 +'1';
		 Energy_Bin_Rdy_1 <= '1';
		else
		 s_Energy_Bin_1 <= s_Energy_Bin_1;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1;   
  
  Energy_Bin_2 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_2   <=  (others =>'0');
	    Energy_Bin_Rdy_2 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E2_C1_L and PEAK_C1 <= s_E2_C1_H and Bin_OR = '0') then
         s_Energy_Bin_2 <= s_Energy_Bin_2 +'1';
		 Energy_Bin_Rdy_2 <= '1';
		else
		 s_Energy_Bin_2 <= s_Energy_Bin_2;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_2 <= '0';
      end if;
    end if;
  end process  Energy_Bin_2;   
  
  Energy_Bin_3 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_3   <=  (others =>'0');
	    Energy_Bin_Rdy_3 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E3_C1_L and PEAK_C1 <= s_E3_C1_H and Bin_OR = '0') then
         s_Energy_Bin_3 <= s_Energy_Bin_3 +'1';
		 Energy_Bin_Rdy_3 <= '1';
		else
		 s_Energy_Bin_3 <= s_Energy_Bin_3;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_3 <= '0';
      end if;
    end if;
  end process  Energy_Bin_3;   
  
  Energy_Bin_4 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_4   <=  (others =>'0');
		Energy_Bin_Rdy_4 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E4_C1_L and PEAK_C1 <= s_E4_C1_H and Bin_OR = '0') then
         s_Energy_Bin_4 <= s_Energy_Bin_4 +'1';
		 Energy_Bin_Rdy_4 <= '1';
		else
		 s_Energy_Bin_4 <= s_Energy_Bin_4;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_4 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_4;   
 
 
  Energy_Bin_5 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_5   <=  (others =>'0');
		Energy_Bin_Rdy_5 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E5_C1_L and PEAK_C1 <= s_E5_C1_H and Bin_OR = '0') then
         s_Energy_Bin_5 <= s_Energy_Bin_5 +'1';
		 Energy_Bin_Rdy_5 <= '1';
		else
		 s_Energy_Bin_5 <= s_Energy_Bin_5;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_5 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_5;  
 
  
  Energy_Bin_6 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_6   <=  (others =>'0');
		Energy_Bin_Rdy_6 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E6_C1_L and PEAK_C1 <= s_E6_C1_H and Bin_OR = '0') then
         s_Energy_Bin_6 <= s_Energy_Bin_6 +'1';
		 Energy_Bin_Rdy_6 <= '1';
		else
		 s_Energy_Bin_6 <= s_Energy_Bin_6;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_6 <= '0';
      end if;
    end if;
  end process  Energy_Bin_6;   
  
 Energy_Bin_7 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_7   <=  (others =>'0');
		Energy_Bin_Rdy_7 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E7_C1_L and PEAK_C1 <= s_E7_C1_H and Bin_OR = '0') then
         s_Energy_Bin_7 <= s_Energy_Bin_7 +'1';
		 Energy_Bin_Rdy_7 <= '1';
		else
		 s_Energy_Bin_7 <= s_Energy_Bin_7;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_7 <= '0';
      end if;
    end if;
  end process  Energy_Bin_7;   
  
  Energy_Bin_8 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_8   <=  (others =>'0');
		Energy_Bin_Rdy_8 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E8_C1_L and PEAK_C1 <= s_E8_C1_H and Bin_OR = '0') then
         s_Energy_Bin_8 <= s_Energy_Bin_8 +'1';
		 Energy_Bin_Rdy_8 <= '1';
		else
		 s_Energy_Bin_8 <= s_Energy_Bin_8;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_8 <= '0';
      end if;
    end if;
  end process  Energy_Bin_8;   
  
  Energy_Bin_9 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_9   <=  (others =>'0');
		Energy_Bin_Rdy_9 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E9_C1_L and PEAK_C1 <= s_E9_C1_H and Bin_OR = '0') then
         s_Energy_Bin_9 <= s_Energy_Bin_9 +'1';
		 Energy_Bin_Rdy_9 <= '1';
		else
		 s_Energy_Bin_9 <= s_Energy_Bin_9;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_9 <= '0';
      end if;
    end if;
  end process  Energy_Bin_9;   
  
  Energy_Bin_10 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_10   <=  (others =>'0');
		Energy_Bin_Rdy_10 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E10_C1_L and PEAK_C1 <= s_E10_C1_H and Bin_OR = '0') then
         s_Energy_Bin_10 <= s_Energy_Bin_10 +'1';
		 Energy_Bin_Rdy_10 <= '1';
		else
		 s_Energy_Bin_10 <= s_Energy_Bin_10;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_10 <= '0';
      end if;
    end if;
  end process  Energy_Bin_10;   
  
  Energy_Bin_11 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_11   <=  (others =>'0');
		Energy_Bin_Rdy_11 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E11_C1_L and PEAK_C1 <= s_E11_C1_H and Bin_OR = '0') then
         s_Energy_Bin_11 <= s_Energy_Bin_11 +'1';
		 Energy_Bin_Rdy_11 <= '1';
		else
		 s_Energy_Bin_11 <= s_Energy_Bin_11;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_11 <= '0';
      end if;
    end if;
  end process  Energy_Bin_11;   
  
    Energy_Bin_12 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_12   <=  (others =>'0');
		Energy_Bin_Rdy_12 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E12_C1_L and PEAK_C1 <= s_E12_C1_H and Bin_OR = '0') then
         s_Energy_Bin_12 <= s_Energy_Bin_12 +'1';
		 Energy_Bin_Rdy_12 <= '1';
		else
		 s_Energy_Bin_12 <= s_Energy_Bin_12;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_12 <= '0';
      end if;
    end if;
  end process  Energy_Bin_12;   

    Energy_Bin_13 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_13   <=  (others =>'0');
		Energy_Bin_Rdy_13 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E13_C1_L and PEAK_C1 <= s_E13_C1_H and Bin_OR = '0') then
         s_Energy_Bin_13 <= s_Energy_Bin_13 +'1';
		 Energy_Bin_Rdy_13 <= '1';
		else
		 s_Energy_Bin_13 <= s_Energy_Bin_13;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_13 <= '0';
      end if;
    end if;
  end process  Energy_Bin_13;   
  
     Energy_Bin_14 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_14   <=  (others =>'0');
		Energy_Bin_Rdy_14 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E14_C1_L and PEAK_C1 <= s_E14_C1_H and Bin_OR = '0') then
         s_Energy_Bin_14 <= s_Energy_Bin_14 +'1';
		 Energy_Bin_Rdy_14 <= '1';
		else
		 s_Energy_Bin_14 <= s_Energy_Bin_14;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_14 <= '0';
      end if;
    end if;
  end process  Energy_Bin_14;    
  
     Energy_Bin_15 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_15   <=  (others =>'0');
		Energy_Bin_Rdy_15 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E15_C1_L and PEAK_C1 <= s_E15_C1_H and Bin_OR = '0') then
         s_Energy_Bin_15 <= s_Energy_Bin_15 +'1';
		 Energy_Bin_Rdy_15 <= '1';
		else
		 s_Energy_Bin_15 <= s_Energy_Bin_15;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_15 <= '0';
      end if;
    end if;
  end process  Energy_Bin_15;      
  
     Energy_Bin_16 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_16   <=  (others =>'0');
		Energy_Bin_Rdy_16 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E16_C1_L and PEAK_C1 <= s_E16_C1_H and Bin_OR = '0') then
         s_Energy_Bin_16 <= s_Energy_Bin_16 +'1';
		 Energy_Bin_Rdy_16 <= '1';
		else
		 s_Energy_Bin_16 <= s_Energy_Bin_16;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_16 <= '0';
      end if;
    end if;
  end process  Energy_Bin_16;     
  
     Energy_Bin_17 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_17   <=  (others =>'0');
		Energy_Bin_Rdy_17 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E17_C1_L and PEAK_C1 <= s_E17_C1_H and Bin_OR = '0') then
         s_Energy_Bin_17 <= s_Energy_Bin_17 +'1';
		 Energy_Bin_Rdy_17 <= '1';
		else
		 s_Energy_Bin_17 <= s_Energy_Bin_17;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_17 <= '0';
      end if;
    end if;
  end process  Energy_Bin_17;     
  
     Energy_Bin_18 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_18   <=  (others =>'0');
		Energy_Bin_Rdy_18 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E18_C1_L and PEAK_C1 <= s_E18_C1_H and Bin_OR = '0') then
         s_Energy_Bin_18 <= s_Energy_Bin_18 +'1';
		 Energy_Bin_Rdy_18 <= '1';
		else
		 s_Energy_Bin_18 <= s_Energy_Bin_18;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_18 <= '0';
      end if;
    end if;
  end process  Energy_Bin_18;       
  
     Energy_Bin_19 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_19   <=  (others =>'0');
		Energy_Bin_Rdy_19 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E19_C1_L and PEAK_C1 <= s_E19_C1_H and Bin_OR = '0') then
         s_Energy_Bin_19 <= s_Energy_Bin_19 +'1';
		 Energy_Bin_Rdy_19 <= '1';
		else
		 s_Energy_Bin_19 <= s_Energy_Bin_19;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_19 <= '0';
      end if;
    end if;
  end process  Energy_Bin_19;     
  
      Energy_Bin_20 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_20   <=  (others =>'0');
		Energy_Bin_Rdy_20 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E20_C1_L and PEAK_C1 <= s_E20_C1_H and Bin_OR = '0') then
         s_Energy_Bin_20 <= s_Energy_Bin_20 +'1';
		 Energy_Bin_Rdy_20 <= '1';
		else
		 s_Energy_Bin_20 <= s_Energy_Bin_20;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_20 <= '0';
      end if;
    end if;
  end process  Energy_Bin_20;      
  
  Energy_Bin_21 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_21   <=  (others =>'0');
		Energy_Bin_Rdy_21 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E21_C1_L and PEAK_C1 <= s_E21_C1_H and Bin_OR = '0') then
         s_Energy_Bin_21 <= s_Energy_Bin_21 +'1';
		 Energy_Bin_Rdy_21 <= '1';
		else
		 s_Energy_Bin_21 <= s_Energy_Bin_21;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_21 <= '0';
      end if;
    end if;
  end process  Energy_Bin_21;   
  
    Energy_Bin_22 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_22   <=  (others =>'0');
		Energy_Bin_Rdy_22 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E22_C1_L and PEAK_C1 <= s_E22_C1_H and Bin_OR = '0') then
         s_Energy_Bin_22 <= s_Energy_Bin_22 +'1';
		 Energy_Bin_Rdy_22 <= '1';
		else
		 s_Energy_Bin_22 <= s_Energy_Bin_22;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_22 <= '0';
      end if;
    end if;
  end process  Energy_Bin_22;   

    Energy_Bin_23 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_23   <=  (others =>'0');
		Energy_Bin_Rdy_23 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E23_C1_L and PEAK_C1 <= s_E23_C1_H and Bin_OR = '0') then
         s_Energy_Bin_23 <= s_Energy_Bin_23 +'1';
		 Energy_Bin_Rdy_23 <= '1';
		else
		 s_Energy_Bin_23 <= s_Energy_Bin_23;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_23 <= '0';
      end if;
    end if;
  end process  Energy_Bin_23;   
  
     Energy_Bin_24 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_24   <=  (others =>'0');
		Energy_Bin_Rdy_24 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E24_C1_L and PEAK_C1 <= s_E24_C1_H and Bin_OR = '0') then
         s_Energy_Bin_24 <= s_Energy_Bin_24 +'1';
		 Energy_Bin_Rdy_24 <= '1';
		else
		 s_Energy_Bin_24 <= s_Energy_Bin_24;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_24 <= '0';
      end if;
    end if;
  end process  Energy_Bin_24;    
  
     Energy_Bin_25 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_25   <=  (others =>'0');
		Energy_Bin_Rdy_25 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E25_C1_L and PEAK_C1 <= s_E25_C1_H and Bin_OR = '0') then
         s_Energy_Bin_25 <= s_Energy_Bin_25 +'1';
		 Energy_Bin_Rdy_25 <= '1';
		else
		 s_Energy_Bin_25 <= s_Energy_Bin_25;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_25 <= '0';
      end if;
    end if;
  end process  Energy_Bin_25;      
  
     Energy_Bin_26 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_26   <=  (others =>'0');
		Energy_Bin_Rdy_26 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E26_C1_L and PEAK_C1 <= s_E26_C1_H and Bin_OR = '0') then
         s_Energy_Bin_26 <= s_Energy_Bin_26 +'1';
		 Energy_Bin_Rdy_26 <= '1';
		else
		 s_Energy_Bin_26 <= s_Energy_Bin_26;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_26 <= '0';
      end if;
    end if;
  end process  Energy_Bin_26;     
  
     Energy_Bin_27 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_27   <=  (others =>'0');
		Energy_Bin_Rdy_27 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E27_C1_L and PEAK_C1 <= s_E27_C1_H and Bin_OR = '0') then
         s_Energy_Bin_27 <= s_Energy_Bin_27 +'1';
		 Energy_Bin_Rdy_27 <= '1';
		else
		 s_Energy_Bin_27 <= s_Energy_Bin_27;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_27 <= '0';
      end if;
    end if;
  end process  Energy_Bin_27;     
  
     Energy_Bin_28 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_28   <=  (others =>'0');
		Energy_Bin_Rdy_28 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E28_C1_L and PEAK_C1 <= s_E28_C1_H and Bin_OR = '0') then
         s_Energy_Bin_28 <= s_Energy_Bin_28 +'1';
		 Energy_Bin_Rdy_28 <= '1';
		else
		 s_Energy_Bin_28 <= s_Energy_Bin_28;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_28 <= '0';
      end if;
    end if;
  end process  Energy_Bin_28;       
  
     Energy_Bin_29 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_29   <=  (others =>'0');
		Energy_Bin_Rdy_29 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E29_C1_L and PEAK_C1 <= s_E29_C1_H and Bin_OR = '0') then
         s_Energy_Bin_29 <= s_Energy_Bin_29 +'1';
		 Energy_Bin_Rdy_29 <= '1';
		else
		 s_Energy_Bin_29 <= s_Energy_Bin_29;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_29 <= '0';
      end if;
    end if;
  end process  Energy_Bin_29;   

  Energy_Bin_30 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_30   <=  (others =>'0');
		Energy_Bin_Rdy_30 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E30_C1_L and PEAK_C1 <= s_E30_C1_H and Bin_OR = '0') then
         s_Energy_Bin_30 <= s_Energy_Bin_30 +'1';
		 Energy_Bin_Rdy_30 <= '1';
		else
		 s_Energy_Bin_30 <= s_Energy_Bin_30;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_30 <= '0';
      end if;
    end if;
  end process  Energy_Bin_30;     
  
  Energy_Bin_31 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_31   <=  (others =>'0');
		Energy_Bin_Rdy_31 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E31_C1_L and PEAK_C1 <= s_E31_C1_H and Bin_OR = '0') then
         s_Energy_Bin_31 <= s_Energy_Bin_31 +'1';
		 Energy_Bin_Rdy_31 <= '1';
		else
		 s_Energy_Bin_31 <= s_Energy_Bin_31;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_31 <= '0';
      end if;
    end if;
  end process  Energy_Bin_31;   
  
    Energy_Bin_32 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_32   <=  (others =>'0');
		Energy_Bin_Rdy_32 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E32_C1_L and PEAK_C1 <= s_E32_C1_H and Bin_OR = '0') then
         s_Energy_Bin_32 <= s_Energy_Bin_32 +'1';
		 Energy_Bin_Rdy_32 <= '1';
		else
		 s_Energy_Bin_32 <= s_Energy_Bin_32;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_32 <= '0';
      end if;
    end if;
  end process  Energy_Bin_32;   

    Energy_Bin_33 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_33   <=  (others =>'0');
		Energy_Bin_Rdy_33 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E33_C1_L and PEAK_C1 <= s_E33_C1_H and Bin_OR = '0') then
         s_Energy_Bin_33 <= s_Energy_Bin_33 +'1';
		 Energy_Bin_Rdy_33 <= '1';
		else
		 s_Energy_Bin_33 <= s_Energy_Bin_33;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_33 <= '0';
      end if;
    end if;
  end process  Energy_Bin_33;   
  
     Energy_Bin_34 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_34   <=  (others =>'0');
		Energy_Bin_Rdy_34 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E34_C1_L and PEAK_C1 <= s_E34_C1_H and Bin_OR = '0') then
         s_Energy_Bin_34 <= s_Energy_Bin_34 +'1';
		 Energy_Bin_Rdy_34 <= '1';
		else
		 s_Energy_Bin_34 <= s_Energy_Bin_34;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_34 <= '0';
      end if;
    end if;
  end process  Energy_Bin_34;    
  
     Energy_Bin_35 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_35   <=  (others =>'0');
		Energy_Bin_Rdy_35 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E35_C1_L and PEAK_C1 <= s_E35_C1_H and Bin_OR = '0') then
         s_Energy_Bin_35 <= s_Energy_Bin_35 +'1';
		 Energy_Bin_Rdy_35 <= '1';
		else
		 s_Energy_Bin_35 <= s_Energy_Bin_35;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_35 <= '0';
      end if;
    end if;
  end process  Energy_Bin_35;      
  
     Energy_Bin_36 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_36   <=  (others =>'0');
		Energy_Bin_Rdy_36 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E36_C1_L and PEAK_C1 <= s_E36_C1_H and Bin_OR = '0') then
         s_Energy_Bin_36 <= s_Energy_Bin_36 +'1';
		 Energy_Bin_Rdy_36 <= '1';
		else
		 s_Energy_Bin_36 <= s_Energy_Bin_36;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_36 <= '0';
      end if;
    end if;
  end process  Energy_Bin_36;     
  
     Energy_Bin_37 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_37   <=  (others =>'0');
		Energy_Bin_Rdy_37 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E37_C1_L and PEAK_C1 <= s_E37_C1_H and Bin_OR = '0') then
         s_Energy_Bin_37 <= s_Energy_Bin_37 +'1';
		 Energy_Bin_Rdy_37 <= '1';
		else
		 s_Energy_Bin_37 <= s_Energy_Bin_37;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_37 <= '0';
      end if;
    end if;
  end process  Energy_Bin_37;     
  
     Energy_Bin_38 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_38   <=  (others =>'0');
		Energy_Bin_Rdy_38 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E38_C1_L and PEAK_C1 <= s_E38_C1_H and Bin_OR = '0') then
         s_Energy_Bin_38 <= s_Energy_Bin_38 +'1';
		 Energy_Bin_Rdy_38 <= '1';
		else
		 s_Energy_Bin_38 <= s_Energy_Bin_38;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_38 <= '0';
      end if;
    end if;
  end process  Energy_Bin_38;       
  
     Energy_Bin_39 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_39   <=  (others =>'0');
		Energy_Bin_Rdy_39 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E39_C1_L and PEAK_C1 <= s_E39_C1_H and Bin_OR = '0') then
         s_Energy_Bin_39 <= s_Energy_Bin_39 +'1';
		 Energy_Bin_Rdy_39 <= '1';
		else
		 s_Energy_Bin_39 <= s_Energy_Bin_39;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_39 <= '0';
      end if;
    end if;
  end process  Energy_Bin_39;       

  Energy_Bin_40 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_40   <=  (others =>'0');
		Energy_Bin_Rdy_40 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E40_C1_L and PEAK_C1 <= s_E40_C1_H and Bin_OR = '0') then
         s_Energy_Bin_40 <= s_Energy_Bin_40 +'1';
		 Energy_Bin_Rdy_40 <= '1';
		else
		 s_Energy_Bin_40 <= s_Energy_Bin_40;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_40 <= '0';
      end if;
    end if;
  end process  Energy_Bin_40;   
  
  Energy_Bin_41 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_41   <=  (others =>'0');
		Energy_Bin_Rdy_41 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E41_C1_L and PEAK_C1 <= s_E41_C1_H and Bin_OR = '0') then
         s_Energy_Bin_41 <= s_Energy_Bin_41 +'1';
		 Energy_Bin_Rdy_41 <= '1';
		else
		 s_Energy_Bin_41 <= s_Energy_Bin_41;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_41 <= '0';
      end if;
    end if;
  end process  Energy_Bin_41;   
  
    Energy_Bin_42 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_42   <=  (others =>'0');
		Energy_Bin_Rdy_42 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E42_C1_L and PEAK_C1 <= s_E42_C1_H and Bin_OR = '0') then
         s_Energy_Bin_42 <= s_Energy_Bin_42 +'1';
		 Energy_Bin_Rdy_42 <= '1';
		else
		 s_Energy_Bin_42 <= s_Energy_Bin_42;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_42 <= '0';
      end if;
    end if;
  end process  Energy_Bin_42;   

    Energy_Bin_43 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_43   <=  (others =>'0');
		Energy_Bin_Rdy_43 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E43_C1_L and PEAK_C1 <= s_E43_C1_H and Bin_OR = '0') then
         s_Energy_Bin_43 <= s_Energy_Bin_43 +'1';
		 Energy_Bin_Rdy_43 <= '1';
		else
		 s_Energy_Bin_43 <= s_Energy_Bin_43;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_43 <= '0';
      end if;
    end if;
  end process  Energy_Bin_43;   
  
     Energy_Bin_44 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_44   <=  (others =>'0');
		Energy_Bin_Rdy_44 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E44_C1_L and PEAK_C1 <= s_E44_C1_H and Bin_OR = '0') then
         s_Energy_Bin_44 <= s_Energy_Bin_44 +'1';
		 Energy_Bin_Rdy_44 <= '1';
		else
		 s_Energy_Bin_44 <= s_Energy_Bin_44;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_44 <= '0';
      end if;
    end if;
  end process  Energy_Bin_44;    
  
     Energy_Bin_45 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_45   <=  (others =>'0');
		Energy_Bin_Rdy_45 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E45_C1_L and PEAK_C1 <= s_E45_C1_H and Bin_OR = '0') then
         s_Energy_Bin_45 <= s_Energy_Bin_45 +'1';
		 Energy_Bin_Rdy_45 <= '1';
		else
		 s_Energy_Bin_45 <= s_Energy_Bin_45;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_45 <= '0';
      end if;
    end if;
  end process  Energy_Bin_45;      
  
     Energy_Bin_46 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_46   <=  (others =>'0');
		Energy_Bin_Rdy_46 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E46_C1_L and PEAK_C1 <= s_E46_C1_H and Bin_OR = '0') then
         s_Energy_Bin_46 <= s_Energy_Bin_46 +'1';
		 Energy_Bin_Rdy_46 <= '1';
		else
		 s_Energy_Bin_46 <= s_Energy_Bin_46;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_46 <= '0';
      end if;
    end if;
  end process  Energy_Bin_46;     
  
     Energy_Bin_47 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_47   <=  (others =>'0');
		Energy_Bin_Rdy_47 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E47_C1_L and PEAK_C1 <= s_E47_C1_H and Bin_OR = '0') then
         s_Energy_Bin_47 <= s_Energy_Bin_47 +'1';
		 Energy_Bin_Rdy_47 <= '1';
		else
		 s_Energy_Bin_47 <= s_Energy_Bin_47;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_47 <= '0';
      end if;
    end if;
  end process  Energy_Bin_47;     
  
     Energy_Bin_48 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_48   <=  (others =>'0');
		Energy_Bin_Rdy_48 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E48_C1_L and PEAK_C1 <= s_E48_C1_H and Bin_OR = '0') then
         s_Energy_Bin_48 <= s_Energy_Bin_48 +'1';
		 Energy_Bin_Rdy_48 <= '1';
		else
		 s_Energy_Bin_48 <= s_Energy_Bin_48;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_48 <= '0';
      end if;
    end if;
  end process  Energy_Bin_48;       
  
     Energy_Bin_49 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_49   <=  (others =>'0');
		Energy_Bin_Rdy_49 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E49_C1_L and PEAK_C1 <= s_E49_C1_H and Bin_OR = '0') then
         s_Energy_Bin_49 <= s_Energy_Bin_49 +'1';
		 Energy_Bin_Rdy_49 <= '1';
		else
		 s_Energy_Bin_49 <= s_Energy_Bin_49;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_49 <= '0';
      end if;
    end if;
  end process  Energy_Bin_49;        
 
  Energy_Bin_50 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_50   <=  (others =>'0');
		Energy_Bin_Rdy_50 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E50_C1_L and PEAK_C1 <= s_E50_C1_H and Bin_OR = '0') then
         s_Energy_Bin_50 <= s_Energy_Bin_50 +'1';
		 Energy_Bin_Rdy_50 <= '1';
		else
		 s_Energy_Bin_50 <= s_Energy_Bin_50;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_50 <= '0';
      end if;
    end if;
  end process  Energy_Bin_50;   
  
  Energy_Bin_51 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_51   <=  (others =>'0');
		Energy_Bin_Rdy_51 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E51_C1_L and PEAK_C1 <= s_E51_C1_H and Bin_OR = '0') then
         s_Energy_Bin_51 <= s_Energy_Bin_51 +'1';
		 Energy_Bin_Rdy_51 <= '1';
		else
		 s_Energy_Bin_51 <= s_Energy_Bin_51;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_51 <= '0';
      end if;
    end if;
  end process  Energy_Bin_51;   
  
    Energy_Bin_52 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_52   <=  (others =>'0');
		Energy_Bin_Rdy_52 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E52_C1_L and PEAK_C1 <= s_E52_C1_H and Bin_OR = '0') then
         s_Energy_Bin_52 <= s_Energy_Bin_52 +'1';
		 Energy_Bin_Rdy_52 <= '1';
		else
		 s_Energy_Bin_52 <= s_Energy_Bin_52;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_52 <= '0';
      end if;
    end if;
  end process  Energy_Bin_52;   

    Energy_Bin_53 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_53   <=  (others =>'0');
		Energy_Bin_Rdy_53 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E53_C1_L and PEAK_C1 <= s_E53_C1_H and Bin_OR = '0') then
         s_Energy_Bin_53 <= s_Energy_Bin_53 +'1';
		 Energy_Bin_Rdy_53 <= '1';
		else
		 s_Energy_Bin_53 <= s_Energy_Bin_53;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_53 <= '0';
      end if;
    end if;
  end process  Energy_Bin_53;   
  
     Energy_Bin_54 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_54   <=  (others =>'0');
		Energy_Bin_Rdy_54 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E54_C1_L and PEAK_C1 <= s_E54_C1_H and Bin_OR = '0') then
         s_Energy_Bin_54 <= s_Energy_Bin_54 +'1';
		 Energy_Bin_Rdy_54 <= '1';
		else
		 s_Energy_Bin_54 <= s_Energy_Bin_54;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_54 <= '0';
      end if;
    end if;
  end process  Energy_Bin_54;    
  
     Energy_Bin_55 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_55   <=  (others =>'0');
		Energy_Bin_Rdy_55 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E55_C1_L and PEAK_C1 <= s_E55_C1_H and Bin_OR = '0') then
         s_Energy_Bin_55 <= s_Energy_Bin_55 +'1';
		 Energy_Bin_Rdy_55 <= '1';
		else
		 s_Energy_Bin_55 <= s_Energy_Bin_55;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_55 <= '0';
      end if;
    end if;
  end process  Energy_Bin_55;      
  
     Energy_Bin_56 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_56   <=  (others =>'0');
		Energy_Bin_Rdy_56 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E56_C1_L and PEAK_C1 <= s_E56_C1_H and Bin_OR = '0') then
         s_Energy_Bin_56 <= s_Energy_Bin_56 +'1';
		 Energy_Bin_Rdy_56 <= '1';
		else
		 s_Energy_Bin_56 <= s_Energy_Bin_56;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_56 <= '0';
      end if;
    end if;
  end process  Energy_Bin_56;     
  
     Energy_Bin_57 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_57   <=  (others =>'0');
		Energy_Bin_Rdy_57 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E57_C1_L and PEAK_C1 <= s_E57_C1_H and Bin_OR = '0') then
         s_Energy_Bin_57 <= s_Energy_Bin_57 +'1';
		 Energy_Bin_Rdy_57 <= '1';
		else
		 s_Energy_Bin_57 <= s_Energy_Bin_57;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_57 <= '0';
      end if;
    end if;
  end process  Energy_Bin_57;     
  
     Energy_Bin_58 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_58   <=  (others =>'0');
		Energy_Bin_Rdy_58 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E58_C1_L and PEAK_C1 <= s_E58_C1_H and Bin_OR = '0') then
         s_Energy_Bin_58 <= s_Energy_Bin_58 +'1';
		 Energy_Bin_Rdy_58 <= '1';
		else
		 s_Energy_Bin_58 <= s_Energy_Bin_58;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_58 <= '0';
      end if;
    end if;
  end process  Energy_Bin_58;       
  
     Energy_Bin_59 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_59   <=  (others =>'0');
		Energy_Bin_Rdy_59 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E59_C1_L and PEAK_C1 <= s_E59_C1_H and Bin_OR = '0') then
         s_Energy_Bin_59 <= s_Energy_Bin_59 +'1';
		 Energy_Bin_Rdy_59 <= '1';
		else
		 s_Energy_Bin_59 <= s_Energy_Bin_59;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_59 <= '0';
      end if;
    end if;
  end process  Energy_Bin_59;        

     Energy_Bin_60 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_60   <=  (others =>'0');
		Energy_Bin_Rdy_60 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E60_C1_L and PEAK_C1 <= s_E60_C1_H and Bin_OR = '0') then
         s_Energy_Bin_60 <= s_Energy_Bin_60 +'1';
		 Energy_Bin_Rdy_60 <= '1';
		else
		 s_Energy_Bin_60 <= s_Energy_Bin_60;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_60 <= '0';
      end if;
    end if;
  end process  Energy_Bin_60; 
  
  Energy_Bin_61 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_61   <=  (others =>'0');
		Energy_Bin_Rdy_61 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E61_C1_L and PEAK_C1 <= s_E61_C1_H and Bin_OR = '0') then
         s_Energy_Bin_61 <= s_Energy_Bin_61 +'1';
		 Energy_Bin_Rdy_61 <= '1';
		else
		 s_Energy_Bin_61 <= s_Energy_Bin_61;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_61 <= '0';
      end if;
    end if;
  end process  Energy_Bin_61;   
  
    Energy_Bin_62 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_62   <=  (others =>'0');
		Energy_Bin_Rdy_62 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E62_C1_L and PEAK_C1 <= s_E62_C1_H and Bin_OR = '0') then
         s_Energy_Bin_62 <= s_Energy_Bin_62 +'1';
		 Energy_Bin_Rdy_62 <= '1';
		else
		 s_Energy_Bin_62 <= s_Energy_Bin_62;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_62 <= '0';
      end if;
    end if;
  end process  Energy_Bin_62;   

    Energy_Bin_63 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_63   <=  (others =>'0');
		Energy_Bin_Rdy_63 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E63_C1_L and PEAK_C1 <= s_E63_C1_H and Bin_OR = '0') then
         s_Energy_Bin_63 <= s_Energy_Bin_63 +'1';
		 Energy_Bin_Rdy_63 <= '1';
		else
		 s_Energy_Bin_63 <= s_Energy_Bin_63;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_63 <= '0';
      end if;
    end if;
  end process  Energy_Bin_63;   
  
     Energy_Bin_64 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_64   <=  (others =>'0');
		Energy_Bin_Rdy_64 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E64_C1_L and PEAK_C1 <= s_E64_C1_H and Bin_OR = '0') then
         s_Energy_Bin_64 <= s_Energy_Bin_64 +'1';
		 Energy_Bin_Rdy_64 <= '1';
		else
		 s_Energy_Bin_64 <= s_Energy_Bin_64;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_64 <= '0';
      end if;
    end if;
  end process  Energy_Bin_64;    
  
     Energy_Bin_65 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_65   <=  (others =>'0');
		Energy_Bin_Rdy_65 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E65_C1_L and PEAK_C1 <= s_E65_C1_H and Bin_OR = '0') then
         s_Energy_Bin_65 <= s_Energy_Bin_65 +'1';
		 Energy_Bin_Rdy_65 <= '1';
		else
		 s_Energy_Bin_65 <= s_Energy_Bin_65;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_65 <= '0';
      end if;
    end if;
  end process  Energy_Bin_65;      
  
     Energy_Bin_66 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_66   <=  (others =>'0');
		Energy_Bin_Rdy_66 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E66_C1_L and PEAK_C1 <= s_E66_C1_H and Bin_OR = '0') then
         s_Energy_Bin_66 <= s_Energy_Bin_66 +'1';
		 Energy_Bin_Rdy_66 <= '1';
		else
		 s_Energy_Bin_66 <= s_Energy_Bin_66;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_66 <= '0';
      end if;
    end if;
  end process  Energy_Bin_66;     
  
     Energy_Bin_67 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_67   <=  (others =>'0');
		Energy_Bin_Rdy_67 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E67_C1_L and PEAK_C1 <= s_E67_C1_H and Bin_OR = '0') then
         s_Energy_Bin_67 <= s_Energy_Bin_67 +'1';
		 Energy_Bin_Rdy_67 <= '1';
		else
		 s_Energy_Bin_67 <= s_Energy_Bin_67;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_67 <= '0';
      end if;
    end if;
  end process  Energy_Bin_67;     
  
     Energy_Bin_68 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_68   <=  (others =>'0');
		Energy_Bin_Rdy_68 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E68_C1_L and PEAK_C1 <= s_E68_C1_H and Bin_OR = '0') then
         s_Energy_Bin_68 <= s_Energy_Bin_68 +'1';
		 Energy_Bin_Rdy_68 <= '1';
		else
		 s_Energy_Bin_68 <= s_Energy_Bin_68;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_68 <= '0';
      end if;
    end if;
  end process  Energy_Bin_68;       
  
     Energy_Bin_69 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_69   <=  (others =>'0');
		Energy_Bin_Rdy_69 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E69_C1_L and PEAK_C1 <= s_E69_C1_H and Bin_OR = '0') then
         s_Energy_Bin_69 <= s_Energy_Bin_69 +'1';
		 Energy_Bin_Rdy_69 <= '1';
		else
		 s_Energy_Bin_69 <= s_Energy_Bin_69;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_69 <= '0';
      end if;
    end if;
  end process  Energy_Bin_69;      

     Energy_Bin_70 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_70   <=  (others =>'0');
		Energy_Bin_Rdy_70 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E70_C1_L and PEAK_C1 <= s_E70_C1_H and Bin_OR = '0') then
         s_Energy_Bin_70 <= s_Energy_Bin_70 +'1';
		 Energy_Bin_Rdy_70 <= '1';
		else
		 s_Energy_Bin_70 <= s_Energy_Bin_70;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_70 <= '0';
      end if;
    end if;
  end process  Energy_Bin_70;       
  
  Energy_Bin_71 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_71   <=  (others =>'0');
		Energy_Bin_Rdy_71 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E71_C1_L and PEAK_C1 <= s_E71_C1_H and Bin_OR = '0') then
         s_Energy_Bin_71 <= s_Energy_Bin_71 +'1';
		 Energy_Bin_Rdy_71 <= '1';
		else
		 s_Energy_Bin_71 <= s_Energy_Bin_71;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_71 <= '0';
      end if;
    end if;
  end process  Energy_Bin_71;   
  
    Energy_Bin_72 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_72   <=  (others =>'0');
		Energy_Bin_Rdy_72 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E72_C1_L and PEAK_C1 <= s_E72_C1_H and Bin_OR = '0') then
         s_Energy_Bin_72 <= s_Energy_Bin_72 +'1';
		 Energy_Bin_Rdy_72 <= '1';
		else
		 s_Energy_Bin_72 <= s_Energy_Bin_72;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_72 <= '0';
      end if;
    end if;
  end process  Energy_Bin_72;   

    Energy_Bin_73 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_73   <=  (others =>'0');
		Energy_Bin_Rdy_73 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E73_C1_L and PEAK_C1 <= s_E73_C1_H and Bin_OR = '0') then
         s_Energy_Bin_73 <= s_Energy_Bin_73 +'1';
		 Energy_Bin_Rdy_73 <= '1';
		else
		 s_Energy_Bin_73 <= s_Energy_Bin_73;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_73 <= '0';
      end if;
    end if;
  end process  Energy_Bin_73;   
  
     Energy_Bin_74 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_74   <=  (others =>'0');
		Energy_Bin_Rdy_74 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E74_C1_L and PEAK_C1 <= s_E74_C1_H and Bin_OR = '0') then
         s_Energy_Bin_74 <= s_Energy_Bin_74 +'1';
		 Energy_Bin_Rdy_74 <= '1';
		else
		 s_Energy_Bin_74 <= s_Energy_Bin_74;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_74 <= '0';
      end if;
    end if;
  end process  Energy_Bin_74;    
  
     Energy_Bin_75 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_75   <=  (others =>'0');
		Energy_Bin_Rdy_75 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E75_C1_L and PEAK_C1 <= s_E75_C1_H and Bin_OR = '0') then
         s_Energy_Bin_75 <= s_Energy_Bin_75 +'1';
		 Energy_Bin_Rdy_75 <= '1';
		else
		 s_Energy_Bin_75 <= s_Energy_Bin_75;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_75 <= '0';
      end if;
    end if;
  end process  Energy_Bin_75;      
  
     Energy_Bin_76 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_76   <=  (others =>'0');
		Energy_Bin_Rdy_76 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E76_C1_L and PEAK_C1 <= s_E76_C1_H and Bin_OR = '0') then
         s_Energy_Bin_76 <= s_Energy_Bin_76 +'1';
		 Energy_Bin_Rdy_76 <= '1';
		else
		 s_Energy_Bin_76 <= s_Energy_Bin_76;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_76 <= '0';
      end if;
    end if;
  end process  Energy_Bin_76;     
  
     Energy_Bin_77 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_77   <=  (others =>'0');
		Energy_Bin_Rdy_77 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E77_C1_L and PEAK_C1 <= s_E77_C1_H and Bin_OR = '0') then
         s_Energy_Bin_77 <= s_Energy_Bin_77 +'1';
		 Energy_Bin_Rdy_77 <= '1';
		else
		 s_Energy_Bin_77 <= s_Energy_Bin_77;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_77 <= '0';
      end if;
    end if;
  end process  Energy_Bin_77;     
  
     Energy_Bin_78 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_78   <=  (others =>'0');
		Energy_Bin_Rdy_78 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E78_C1_L and PEAK_C1 <= s_E78_C1_H and Bin_OR = '0') then
         s_Energy_Bin_78 <= s_Energy_Bin_78 +'1';
		 Energy_Bin_Rdy_78 <= '1';
		else
		 s_Energy_Bin_78 <= s_Energy_Bin_78;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_78 <= '0';
      end if;
    end if;
  end process  Energy_Bin_78;       
  
     Energy_Bin_79 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_79   <=  (others =>'0');
		Energy_Bin_Rdy_79 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E79_C1_L and PEAK_C1 <= s_E79_C1_H and Bin_OR = '0') then
         s_Energy_Bin_79 <= s_Energy_Bin_79 +'1';
		 Energy_Bin_Rdy_79 <= '1';
		else
		 s_Energy_Bin_79 <= s_Energy_Bin_79;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_79 <= '0';
      end if;
    end if;
  end process  Energy_Bin_79;    
  
     Energy_Bin_80 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_80   <=  (others =>'0');
		Energy_Bin_Rdy_80 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E80_C1_L and PEAK_C1 <= s_E80_C1_H and Bin_OR = '0') then
         s_Energy_Bin_80 <= s_Energy_Bin_80 +'1';
		 Energy_Bin_Rdy_80 <= '1';
		else
		 s_Energy_Bin_80 <= s_Energy_Bin_80;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_80 <= '0';
      end if;
    end if;
  end process  Energy_Bin_80;       
  
  Energy_Bin_81 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_81   <=  (others =>'0');
		Energy_Bin_Rdy_81 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E81_C1_L and PEAK_C1 <= s_E81_C1_H and Bin_OR = '0') then
         s_Energy_Bin_81 <= s_Energy_Bin_81 +'1';
		 Energy_Bin_Rdy_81 <= '1';
		else
		 s_Energy_Bin_81 <= s_Energy_Bin_81;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_81 <= '0';
      end if;
    end if;
  end process  Energy_Bin_81;   
  
    Energy_Bin_82 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_82   <=  (others =>'0');
		Energy_Bin_Rdy_82 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E82_C1_L and PEAK_C1 <= s_E82_C1_H and Bin_OR = '0') then
         s_Energy_Bin_82 <= s_Energy_Bin_82 +'1';
		 Energy_Bin_Rdy_82 <= '1';
		else
		 s_Energy_Bin_82 <= s_Energy_Bin_82;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_82 <= '0';
      end if;
    end if;
  end process  Energy_Bin_82;   

    Energy_Bin_83 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_83   <=  (others =>'0');
		Energy_Bin_Rdy_83 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E83_C1_L and PEAK_C1 <= s_E83_C1_H and Bin_OR = '0') then
         s_Energy_Bin_83 <= s_Energy_Bin_83 +'1';
		 Energy_Bin_Rdy_83 <= '1';
		else
		 s_Energy_Bin_83 <= s_Energy_Bin_83;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_83 <= '0';
      end if;
    end if;
  end process  Energy_Bin_83;   
  
     Energy_Bin_84 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_84   <=  (others =>'0');
		Energy_Bin_Rdy_84 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E84_C1_L and PEAK_C1 <= s_E84_C1_H and Bin_OR = '0') then
         s_Energy_Bin_84 <= s_Energy_Bin_84 +'1';
		 Energy_Bin_Rdy_84 <= '1';
		else
		 s_Energy_Bin_84 <= s_Energy_Bin_84;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_84 <= '0';
      end if;
    end if;
  end process  Energy_Bin_84;    
  
     Energy_Bin_85 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_85   <=  (others =>'0');
		Energy_Bin_Rdy_85 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E85_C1_L and PEAK_C1 <= s_E85_C1_H and Bin_OR = '0') then
         s_Energy_Bin_85 <= s_Energy_Bin_85 +'1';
		 Energy_Bin_Rdy_85 <= '1';
		else
		 s_Energy_Bin_85 <= s_Energy_Bin_85;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_85 <= '0';
      end if;
    end if;
  end process  Energy_Bin_85;      
  
     Energy_Bin_86 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_86   <=  (others =>'0');
		Energy_Bin_Rdy_86 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E86_C1_L and PEAK_C1 <= s_E86_C1_H and Bin_OR = '0') then
         s_Energy_Bin_86 <= s_Energy_Bin_86 +'1';
		 Energy_Bin_Rdy_86 <= '1';
		else
		 s_Energy_Bin_86 <= s_Energy_Bin_86;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_86 <= '0';
      end if;
    end if;
  end process  Energy_Bin_86;     
  
     Energy_Bin_87 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_87   <=  (others =>'0');
		Energy_Bin_Rdy_87 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E87_C1_L and PEAK_C1 <= s_E87_C1_H and Bin_OR = '0') then
         s_Energy_Bin_87 <= s_Energy_Bin_87 +'1';
		 Energy_Bin_Rdy_87 <= '1';
		else
		 s_Energy_Bin_87 <= s_Energy_Bin_87;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_87 <= '0';
      end if;
    end if;
  end process  Energy_Bin_87;     
  
     Energy_Bin_88 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_88   <=  (others =>'0');
		Energy_Bin_Rdy_88 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E88_C1_L and PEAK_C1 <= s_E88_C1_H and Bin_OR = '0') then
         s_Energy_Bin_88 <= s_Energy_Bin_88 +'1';
		 Energy_Bin_Rdy_88 <= '1';
		else
		 s_Energy_Bin_88 <= s_Energy_Bin_88;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_88 <= '0';
      end if;
    end if;
  end process  Energy_Bin_88;       
  
     Energy_Bin_89 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_89   <=  (others =>'0');
		Energy_Bin_Rdy_89 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E89_C1_L and PEAK_C1 <= s_E89_C1_H and Bin_OR = '0') then
         s_Energy_Bin_89 <= s_Energy_Bin_89 +'1';
		 Energy_Bin_Rdy_89 <= '1';
		else
		 s_Energy_Bin_89 <= s_Energy_Bin_89;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_89 <= '0';
      end if;
    end if;
  end process  Energy_Bin_89;      

     Energy_Bin_90 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_90   <=  (others =>'0');
		Energy_Bin_Rdy_90 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E90_C1_L and PEAK_C1 <= s_E90_C1_H and Bin_OR = '0') then
         s_Energy_Bin_90 <= s_Energy_Bin_90 +'1';
		 Energy_Bin_Rdy_90 <= '1';
		else
		 s_Energy_Bin_90 <= s_Energy_Bin_90;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_90 <= '0';
      end if;
    end if;
  end process  Energy_Bin_90;       
  
  Energy_Bin_91 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_91   <=  (others =>'0');
		Energy_Bin_Rdy_91 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E91_C1_L and PEAK_C1 <= s_E91_C1_H and Bin_OR = '0') then
         s_Energy_Bin_91 <= s_Energy_Bin_91 +'1';
		 Energy_Bin_Rdy_91 <= '1';
		else
		 s_Energy_Bin_91 <= s_Energy_Bin_91;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_91 <= '0';
      end if;
    end if;
  end process  Energy_Bin_91;   
  
    Energy_Bin_92 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_92   <=  (others =>'0');
		Energy_Bin_Rdy_92 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E92_C1_L and PEAK_C1 <= s_E92_C1_H and Bin_OR = '0') then
         s_Energy_Bin_92 <= s_Energy_Bin_92 +'1';
		 Energy_Bin_Rdy_92 <= '1';
		else
		 s_Energy_Bin_92 <= s_Energy_Bin_92;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_92 <= '0';
      end if;
    end if;
  end process  Energy_Bin_92;   

    Energy_Bin_93 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_93   <=  (others =>'0');
		Energy_Bin_Rdy_93 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E93_C1_L and PEAK_C1 <= s_E93_C1_H and Bin_OR = '0') then
         s_Energy_Bin_93 <= s_Energy_Bin_93 +'1';
		 Energy_Bin_Rdy_93 <= '1';
		else
		 s_Energy_Bin_93 <= s_Energy_Bin_93;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_93 <= '0';
      end if;
    end if;
  end process  Energy_Bin_93;   
  
     Energy_Bin_94 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_94   <=  (others =>'0');
		Energy_Bin_Rdy_94 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E94_C1_L and PEAK_C1 <= s_E94_C1_H and Bin_OR = '0') then
         s_Energy_Bin_94 <= s_Energy_Bin_94 +'1';
		 Energy_Bin_Rdy_94 <= '1';
		else
		 s_Energy_Bin_94 <= s_Energy_Bin_94;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_94 <= '0';
      end if;
    end if;
  end process  Energy_Bin_94;    
  
     Energy_Bin_95 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_95   <=  (others =>'0');
		Energy_Bin_Rdy_95 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E95_C1_L and PEAK_C1 <= s_E95_C1_H and Bin_OR = '0') then
         s_Energy_Bin_95 <= s_Energy_Bin_95 +'1';
		 Energy_Bin_Rdy_95 <= '1';
		else
		 s_Energy_Bin_95 <= s_Energy_Bin_95;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_95 <= '0';
      end if;
    end if;
  end process  Energy_Bin_95;      
  
     Energy_Bin_96 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_96   <=  (others =>'0');
		Energy_Bin_Rdy_96 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E96_C1_L and PEAK_C1 <= s_E96_C1_H and Bin_OR = '0') then
         s_Energy_Bin_96 <= s_Energy_Bin_96 +'1';
		 Energy_Bin_Rdy_96 <= '1';
		else
		 s_Energy_Bin_96 <= s_Energy_Bin_96;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_96 <= '0';
      end if;
    end if;
  end process  Energy_Bin_96;     
  
     Energy_Bin_97 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_97   <=  (others =>'0');
		Energy_Bin_Rdy_97 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E97_C1_L and PEAK_C1 <= s_E97_C1_H and Bin_OR = '0') then
         s_Energy_Bin_97 <= s_Energy_Bin_97 +'1';
		 Energy_Bin_Rdy_97 <= '1';
		else
		 s_Energy_Bin_97 <= s_Energy_Bin_97;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_97 <= '0';
      end if;
    end if;
  end process  Energy_Bin_97;     
  
     Energy_Bin_98 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_98   <=  (others =>'0');
		Energy_Bin_Rdy_98 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E98_C1_L and PEAK_C1 <= s_E98_C1_H and Bin_OR = '0') then
         s_Energy_Bin_98 <= s_Energy_Bin_98 +'1';
		 Energy_Bin_Rdy_98 <= '1';
		else
		 s_Energy_Bin_98 <= s_Energy_Bin_98;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_98 <= '0';
      end if;
    end if;
  end process  Energy_Bin_98;       
  
     Energy_Bin_99 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_99   <=  (others =>'0');
		Energy_Bin_Rdy_99 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E99_C1_L and PEAK_C1 <= s_E99_C1_H and Bin_OR = '0') then
         s_Energy_Bin_99 <= s_Energy_Bin_99 +'1';
		 Energy_Bin_Rdy_99 <= '1';
		else
		 s_Energy_Bin_99 <= s_Energy_Bin_99;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_99 <= '0';
      end if;
    end if;
  end process  Energy_Bin_99;      
  
     Energy_Bin_100 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_100   <=  (others =>'0');
		Energy_Bin_Rdy_100 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E100_C1_L and PEAK_C1 <= s_E100_C1_H and Bin_OR = '0') then
         s_Energy_Bin_100 <= s_Energy_Bin_100 +'1';
		 Energy_Bin_Rdy_100 <= '1';
		else
		 s_Energy_Bin_100 <= s_Energy_Bin_100;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_100 <= '0';
      end if;
    end if;
  end process  Energy_Bin_100;    
  
  Energy_Bin_101 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_101   <=  (others =>'0');
		Energy_Bin_Rdy_101 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E101_C1_L and PEAK_C1 <= s_E101_C1_H and Bin_OR = '0') then
         s_Energy_Bin_101 <= s_Energy_Bin_101 +'1';
		 Energy_Bin_Rdy_101 <= '1';
		else
		 s_Energy_Bin_101 <= s_Energy_Bin_101;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_101 <= '0';
      end if;
    end if;
  end process  Energy_Bin_101;   
  
  Energy_Bin_102 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_102   <=  (others =>'0');
	    Energy_Bin_Rdy_102 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E102_C1_L and PEAK_C1 <= s_E102_C1_H and Bin_OR = '0') then
         s_Energy_Bin_102 <= s_Energy_Bin_102 +'1';
		 Energy_Bin_Rdy_102 <= '1';
		else
		 s_Energy_Bin_102 <= s_Energy_Bin_102;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_102 <= '0';
      end if;
    end if;
  end process  Energy_Bin_102;   
  
  Energy_Bin_103 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_103   <=  (others =>'0');
	    Energy_Bin_Rdy_103 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E103_C1_L and PEAK_C1 <= s_E103_C1_H and Bin_OR = '0') then
         s_Energy_Bin_103 <= s_Energy_Bin_103 +'1';
		 Energy_Bin_Rdy_103 <= '1';
		else
		 s_Energy_Bin_103 <= s_Energy_Bin_103;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_103 <= '0';
      end if;
    end if;
  end process  Energy_Bin_103;   
  
  Energy_Bin_104 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_104   <=  (others =>'0');
		Energy_Bin_Rdy_104 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E104_C1_L and PEAK_C1 <= s_E104_C1_H and Bin_OR = '0') then
         s_Energy_Bin_104 <= s_Energy_Bin_104 +'1';
		 Energy_Bin_Rdy_104 <= '1';
		else
		 s_Energy_Bin_104 <= s_Energy_Bin_104;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_104 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_104;   
 
 
  Energy_Bin_105 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_105   <=  (others =>'0');
		Energy_Bin_Rdy_105 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E105_C1_L and PEAK_C1 <= s_E105_C1_H and Bin_OR = '0') then
         s_Energy_Bin_105 <= s_Energy_Bin_105 +'1';
		 Energy_Bin_Rdy_105 <= '1';
		else
		 s_Energy_Bin_105 <= s_Energy_Bin_105;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_105 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_105;  
 
  
  Energy_Bin_106 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_106   <=  (others =>'0');
		Energy_Bin_Rdy_106 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E106_C1_L and PEAK_C1 <= s_E106_C1_H and Bin_OR = '0') then
         s_Energy_Bin_106 <= s_Energy_Bin_106 +'1';
		 Energy_Bin_Rdy_106 <= '1';
		else
		 s_Energy_Bin_106 <= s_Energy_Bin_106;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_106 <= '0';
      end if;
    end if;
  end process  Energy_Bin_106;   
  
 Energy_Bin_107 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_107   <=  (others =>'0');
		Energy_Bin_Rdy_107 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E107_C1_L and PEAK_C1 <= s_E107_C1_H and Bin_OR = '0') then
         s_Energy_Bin_107 <= s_Energy_Bin_107 +'1';
		 Energy_Bin_Rdy_107 <= '1';
		else
		 s_Energy_Bin_107 <= s_Energy_Bin_107;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_107 <= '0';
      end if;
    end if;
  end process  Energy_Bin_107;   
  
  Energy_Bin_108 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_108   <=  (others =>'0');
		Energy_Bin_Rdy_108 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E108_C1_L and PEAK_C1 <= s_E108_C1_H and Bin_OR = '0') then
         s_Energy_Bin_108 <= s_Energy_Bin_108 +'1';
		 Energy_Bin_Rdy_108 <= '1';
		else
		 s_Energy_Bin_108 <= s_Energy_Bin_108;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_108 <= '0';
      end if;
    end if;
  end process  Energy_Bin_108;   
  
  Energy_Bin_109 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_109   <=  (others =>'0');
		Energy_Bin_Rdy_109 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E109_C1_L and PEAK_C1 <= s_E109_C1_H and Bin_OR = '0') then
         s_Energy_Bin_109 <= s_Energy_Bin_109 +'1';
		 Energy_Bin_Rdy_109 <= '1';
		else
		 s_Energy_Bin_109 <= s_Energy_Bin_109;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_109 <= '0';
      end if;
    end if;
  end process  Energy_Bin_109;     
  
     Energy_Bin_110 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_110   <=  (others =>'0');
		Energy_Bin_Rdy_110 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E110_C1_L and PEAK_C1 <= s_E110_C1_H and Bin_OR = '0') then
         s_Energy_Bin_110 <= s_Energy_Bin_110 +'1';
		 Energy_Bin_Rdy_110 <= '1';
		else
		 s_Energy_Bin_110 <= s_Energy_Bin_110;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_110 <= '0';
      end if;
    end if;
  end process  Energy_Bin_110;    
  
  Energy_Bin_111 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_111   <=  (others =>'0');
		Energy_Bin_Rdy_111 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E111_C1_L and PEAK_C1 <= s_E111_C1_H and Bin_OR = '0') then
         s_Energy_Bin_111 <= s_Energy_Bin_111 +'1';
		 Energy_Bin_Rdy_111 <= '1';
		else
		 s_Energy_Bin_111 <= s_Energy_Bin_111;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_111 <= '0';
      end if;
    end if;
  end process  Energy_Bin_111;   
  
  Energy_Bin_112 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_112   <=  (others =>'0');
	    Energy_Bin_Rdy_112 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E112_C1_L and PEAK_C1 <= s_E112_C1_H and Bin_OR = '0') then
         s_Energy_Bin_112 <= s_Energy_Bin_112 +'1';
		 Energy_Bin_Rdy_112 <= '1';
		else
		 s_Energy_Bin_112 <= s_Energy_Bin_112;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_112 <= '0';
      end if;
    end if;
  end process  Energy_Bin_112;   
  
  Energy_Bin_113 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_113   <=  (others =>'0');
	    Energy_Bin_Rdy_113 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E113_C1_L and PEAK_C1 <= s_E113_C1_H and Bin_OR = '0') then
         s_Energy_Bin_113 <= s_Energy_Bin_113 +'1';
		 Energy_Bin_Rdy_113 <= '1';
		else
		 s_Energy_Bin_113 <= s_Energy_Bin_113;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_113 <= '0';
      end if;
    end if;
  end process  Energy_Bin_113;   
  
  Energy_Bin_114 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_114   <=  (others =>'0');
		Energy_Bin_Rdy_114 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E114_C1_L and PEAK_C1 <= s_E114_C1_H and Bin_OR = '0') then
         s_Energy_Bin_114 <= s_Energy_Bin_114 +'1';
		 Energy_Bin_Rdy_114 <= '1';
		else
		 s_Energy_Bin_114 <= s_Energy_Bin_114;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_114 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_114;   
 
 
  Energy_Bin_115 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_115   <=  (others =>'0');
		Energy_Bin_Rdy_115 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E115_C1_L and PEAK_C1 <= s_E115_C1_H and Bin_OR = '0') then
         s_Energy_Bin_115 <= s_Energy_Bin_115 +'1';
		 Energy_Bin_Rdy_115 <= '1';
		else
		 s_Energy_Bin_115 <= s_Energy_Bin_115;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_115 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_115;  
 
  
  Energy_Bin_116 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_116   <=  (others =>'0');
		Energy_Bin_Rdy_116 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E116_C1_L and PEAK_C1 <= s_E116_C1_H and Bin_OR = '0') then
         s_Energy_Bin_116 <= s_Energy_Bin_116 +'1';
		 Energy_Bin_Rdy_116 <= '1';
		else
		 s_Energy_Bin_116 <= s_Energy_Bin_116;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_116 <= '0';
      end if;
    end if;
  end process  Energy_Bin_116;   
  
 Energy_Bin_117 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_117   <=  (others =>'0');
		Energy_Bin_Rdy_117 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E117_C1_L and PEAK_C1 <= s_E117_C1_H and Bin_OR = '0') then
         s_Energy_Bin_117 <= s_Energy_Bin_117 +'1';
		 Energy_Bin_Rdy_117 <= '1';
		else
		 s_Energy_Bin_117 <= s_Energy_Bin_117;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_117 <= '0';
      end if;
    end if;
  end process  Energy_Bin_117;   
  
  Energy_Bin_118 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_118   <=  (others =>'0');
		Energy_Bin_Rdy_118 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E118_C1_L and PEAK_C1 <= s_E118_C1_H and Bin_OR = '0') then
         s_Energy_Bin_118 <= s_Energy_Bin_118 +'1';
		 Energy_Bin_Rdy_118 <= '1';
		else
		 s_Energy_Bin_118 <= s_Energy_Bin_118;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_118 <= '0';
      end if;
    end if;
  end process  Energy_Bin_118;   
  
  Energy_Bin_119 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_119   <=  (others =>'0');
		Energy_Bin_Rdy_119 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E119_C1_L and PEAK_C1 <= s_E119_C1_H and Bin_OR = '0') then
         s_Energy_Bin_119 <= s_Energy_Bin_119 +'1';
		 Energy_Bin_Rdy_119 <= '1';
		else
		 s_Energy_Bin_119 <= s_Energy_Bin_119;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_119 <= '0';
      end if;
    end if;
  end process  Energy_Bin_119;      
  
     Energy_Bin_120 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_120   <=  (others =>'0');
		Energy_Bin_Rdy_120 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E120_C1_L and PEAK_C1 <= s_E120_C1_H and Bin_OR = '0') then
         s_Energy_Bin_120 <= s_Energy_Bin_120 +'1';
		 Energy_Bin_Rdy_120 <= '1';
		else
		 s_Energy_Bin_120 <= s_Energy_Bin_120;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_120 <= '0';
      end if;
    end if;
  end process  Energy_Bin_120;    
  
  Energy_Bin_121 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_121   <=  (others =>'0');
		Energy_Bin_Rdy_121 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E121_C1_L and PEAK_C1 <= s_E121_C1_H and Bin_OR = '0') then
         s_Energy_Bin_121 <= s_Energy_Bin_121 +'1';
		 Energy_Bin_Rdy_121 <= '1';
		else
		 s_Energy_Bin_121 <= s_Energy_Bin_121;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_121 <= '0';
      end if;
    end if;
  end process  Energy_Bin_121;   
  
  Energy_Bin_122 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_122   <=  (others =>'0');
	    Energy_Bin_Rdy_122 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E122_C1_L and PEAK_C1 <= s_E122_C1_H and Bin_OR = '0') then
         s_Energy_Bin_122 <= s_Energy_Bin_122 +'1';
		 Energy_Bin_Rdy_122 <= '1';
		else
		 s_Energy_Bin_122 <= s_Energy_Bin_122;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_122 <= '0';
      end if;
    end if;
  end process  Energy_Bin_122;   
  
  Energy_Bin_123 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_123   <=  (others =>'0');
	    Energy_Bin_Rdy_123 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E123_C1_L and PEAK_C1 <= s_E123_C1_H and Bin_OR = '0') then
         s_Energy_Bin_123 <= s_Energy_Bin_123 +'1';
		 Energy_Bin_Rdy_123 <= '1';
		else
		 s_Energy_Bin_123 <= s_Energy_Bin_123;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_123 <= '0';
      end if;
    end if;
  end process  Energy_Bin_123;   
  
  Energy_Bin_124 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_124   <=  (others =>'0');
		Energy_Bin_Rdy_124 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E124_C1_L and PEAK_C1 <= s_E124_C1_H and Bin_OR = '0') then
         s_Energy_Bin_124 <= s_Energy_Bin_124 +'1';
		 Energy_Bin_Rdy_124 <= '1';
		else
		 s_Energy_Bin_124 <= s_Energy_Bin_124;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_124 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_124;   
 
 
  Energy_Bin_125 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_125   <=  (others =>'0');
		Energy_Bin_Rdy_125 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E125_C1_L and PEAK_C1 <= s_E125_C1_H and Bin_OR = '0') then
         s_Energy_Bin_125 <= s_Energy_Bin_125 +'1';
		 Energy_Bin_Rdy_125 <= '1';
		else
		 s_Energy_Bin_125 <= s_Energy_Bin_125;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_125 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_125;  
 
  
  Energy_Bin_126 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_126   <=  (others =>'0');
		Energy_Bin_Rdy_126 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E126_C1_L and PEAK_C1 <= s_E126_C1_H and Bin_OR = '0') then
         s_Energy_Bin_126 <= s_Energy_Bin_126 +'1';
		 Energy_Bin_Rdy_126 <= '1';
		else
		 s_Energy_Bin_126 <= s_Energy_Bin_126;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_126 <= '0';
      end if;
    end if;
  end process  Energy_Bin_126;   
  
 Energy_Bin_127 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_127   <=  (others =>'0');
		Energy_Bin_Rdy_127 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E127_C1_L and PEAK_C1 <= s_E127_C1_H and Bin_OR = '0') then
         s_Energy_Bin_127 <= s_Energy_Bin_127 +'1';
		 Energy_Bin_Rdy_127 <= '1';
		else
		 s_Energy_Bin_127 <= s_Energy_Bin_127;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_127 <= '0';
      end if;
    end if;
  end process  Energy_Bin_127;   
  
  Energy_Bin_128 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_128   <=  (others =>'0');
		Energy_Bin_Rdy_128 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E128_C1_L and PEAK_C1 <= s_E128_C1_H and Bin_OR = '0') then
         s_Energy_Bin_128 <= s_Energy_Bin_128 +'1';
		 Energy_Bin_Rdy_128 <= '1';
		else
		 s_Energy_Bin_128 <= s_Energy_Bin_128;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_128 <= '0';
      end if;
    end if;
  end process  Energy_Bin_128;   
  
  Energy_Bin_129 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_129   <=  (others =>'0');
		Energy_Bin_Rdy_129 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E129_C1_L and PEAK_C1 <= s_E129_C1_H and Bin_OR = '0') then
         s_Energy_Bin_129 <= s_Energy_Bin_129 +'1';
		 Energy_Bin_Rdy_129 <= '1';
		else
		 s_Energy_Bin_129 <= s_Energy_Bin_129;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_129 <= '0';
      end if;
    end if;
  end process  Energy_Bin_129;       
  
     Energy_Bin_130 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_130   <=  (others =>'0');
		Energy_Bin_Rdy_130 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E130_C1_L and PEAK_C1 <= s_E130_C1_H and Bin_OR = '0') then
         s_Energy_Bin_130 <= s_Energy_Bin_130 +'1';
		 Energy_Bin_Rdy_130 <= '1';
		else
		 s_Energy_Bin_130 <= s_Energy_Bin_130;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_130 <= '0';
      end if;
    end if;
  end process  Energy_Bin_130;    
  
  Energy_Bin_131 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_131   <=  (others =>'0');
		Energy_Bin_Rdy_131 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E131_C1_L and PEAK_C1 <= s_E131_C1_H and Bin_OR = '0') then
         s_Energy_Bin_131 <= s_Energy_Bin_131 +'1';
		 Energy_Bin_Rdy_131 <= '1';
		else
		 s_Energy_Bin_131 <= s_Energy_Bin_131;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_131 <= '0';
      end if;
    end if;
  end process  Energy_Bin_131;   
  
  Energy_Bin_132 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_132   <=  (others =>'0');
	    Energy_Bin_Rdy_132 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E132_C1_L and PEAK_C1 <= s_E132_C1_H and Bin_OR = '0') then
         s_Energy_Bin_132 <= s_Energy_Bin_132 +'1';
		 Energy_Bin_Rdy_132 <= '1';
		else
		 s_Energy_Bin_132 <= s_Energy_Bin_132;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_132 <= '0';
      end if;
    end if;
  end process  Energy_Bin_132;   
  
  Energy_Bin_133 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_133   <=  (others =>'0');
	    Energy_Bin_Rdy_133 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E133_C1_L and PEAK_C1 <= s_E133_C1_H and Bin_OR = '0') then
         s_Energy_Bin_133 <= s_Energy_Bin_133 +'1';
		 Energy_Bin_Rdy_133 <= '1';
		else
		 s_Energy_Bin_133 <= s_Energy_Bin_133;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_133 <= '0';
      end if;
    end if;
  end process  Energy_Bin_133;   
  
  Energy_Bin_134 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_134   <=  (others =>'0');
		Energy_Bin_Rdy_134 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E134_C1_L and PEAK_C1 <= s_E134_C1_H and Bin_OR = '0') then
         s_Energy_Bin_134 <= s_Energy_Bin_134 +'1';
		 Energy_Bin_Rdy_134 <= '1';
		else
		 s_Energy_Bin_134 <= s_Energy_Bin_134;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_134 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_134;   
 
 
  Energy_Bin_135 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_135   <=  (others =>'0');
		Energy_Bin_Rdy_135 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E135_C1_L and PEAK_C1 <= s_E135_C1_H and Bin_OR = '0') then
         s_Energy_Bin_135 <= s_Energy_Bin_135 +'1';
		 Energy_Bin_Rdy_135 <= '1';
		else
		 s_Energy_Bin_135 <= s_Energy_Bin_135;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_135 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_135;  
 
  
  Energy_Bin_136 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_136   <=  (others =>'0');
		Energy_Bin_Rdy_136 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E136_C1_L and PEAK_C1 <= s_E136_C1_H and Bin_OR = '0') then
         s_Energy_Bin_136 <= s_Energy_Bin_136 +'1';
		 Energy_Bin_Rdy_136 <= '1';
		else
		 s_Energy_Bin_136 <= s_Energy_Bin_136;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_136 <= '0';
      end if;
    end if;
  end process  Energy_Bin_136;   
  
 Energy_Bin_137 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_137   <=  (others =>'0');
		Energy_Bin_Rdy_137 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E137_C1_L and PEAK_C1 <= s_E137_C1_H and Bin_OR = '0') then
         s_Energy_Bin_137 <= s_Energy_Bin_137 +'1';
		 Energy_Bin_Rdy_137 <= '1';
		else
		 s_Energy_Bin_137 <= s_Energy_Bin_137;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_137 <= '0';
      end if;
    end if;
  end process  Energy_Bin_137;   
  
  Energy_Bin_138 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_138   <=  (others =>'0');
		Energy_Bin_Rdy_138 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E138_C1_L and PEAK_C1 <= s_E138_C1_H and Bin_OR = '0') then
         s_Energy_Bin_138 <= s_Energy_Bin_138 +'1';
		 Energy_Bin_Rdy_138 <= '1';
		else
		 s_Energy_Bin_138 <= s_Energy_Bin_138;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_138 <= '0';
      end if;
    end if;
  end process  Energy_Bin_138;   
  
  Energy_Bin_139 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_139   <=  (others =>'0');
		Energy_Bin_Rdy_139 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E139_C1_L and PEAK_C1 <= s_E139_C1_H and Bin_OR = '0') then
         s_Energy_Bin_139 <= s_Energy_Bin_139 +'1';
		 Energy_Bin_Rdy_139 <= '1';
		else
		 s_Energy_Bin_139 <= s_Energy_Bin_139;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_139 <= '0';
      end if;
    end if;
  end process  Energy_Bin_139;         
  
     Energy_Bin_140 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_140   <=  (others =>'0');
		Energy_Bin_Rdy_140 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E140_C1_L and PEAK_C1 <= s_E140_C1_H and Bin_OR = '0') then
         s_Energy_Bin_140 <= s_Energy_Bin_140 +'1';
		 Energy_Bin_Rdy_140 <= '1';
		else
		 s_Energy_Bin_140 <= s_Energy_Bin_140;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_140 <= '0';
      end if;
    end if;
  end process  Energy_Bin_140;    
  
  Energy_Bin_141 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_141   <=  (others =>'0');
		Energy_Bin_Rdy_141 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E141_C1_L and PEAK_C1 <= s_E141_C1_H and Bin_OR = '0') then
         s_Energy_Bin_141 <= s_Energy_Bin_141 +'1';
		 Energy_Bin_Rdy_141 <= '1';
		else
		 s_Energy_Bin_141 <= s_Energy_Bin_141;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_141 <= '0';
      end if;
    end if;
  end process  Energy_Bin_141;   
  
  Energy_Bin_142 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_142   <=  (others =>'0');
	    Energy_Bin_Rdy_142 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E142_C1_L and PEAK_C1 <= s_E142_C1_H and Bin_OR = '0') then
         s_Energy_Bin_142 <= s_Energy_Bin_142 +'1';
		 Energy_Bin_Rdy_142 <= '1';
		else
		 s_Energy_Bin_142 <= s_Energy_Bin_142;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_142 <= '0';
      end if;
    end if;
  end process  Energy_Bin_142;   
  
  Energy_Bin_143 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_143   <=  (others =>'0');
	    Energy_Bin_Rdy_143 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E143_C1_L and PEAK_C1 <= s_E143_C1_H and Bin_OR = '0') then
         s_Energy_Bin_143 <= s_Energy_Bin_143 +'1';
		 Energy_Bin_Rdy_143 <= '1';
		else
		 s_Energy_Bin_143 <= s_Energy_Bin_143;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_143 <= '0';
      end if;
    end if;
  end process  Energy_Bin_143;   
  
  Energy_Bin_144 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_144   <=  (others =>'0');
		Energy_Bin_Rdy_144 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E144_C1_L and PEAK_C1 <= s_E144_C1_H and Bin_OR = '0') then
         s_Energy_Bin_144 <= s_Energy_Bin_144 +'1';
		 Energy_Bin_Rdy_144 <= '1';
		else
		 s_Energy_Bin_144 <= s_Energy_Bin_144;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_144 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_144;   
 
 
  Energy_Bin_145 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_145   <=  (others =>'0');
		Energy_Bin_Rdy_145 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E145_C1_L and PEAK_C1 <= s_E145_C1_H and Bin_OR = '0') then
         s_Energy_Bin_145 <= s_Energy_Bin_145 +'1';
		 Energy_Bin_Rdy_145 <= '1';
		else
		 s_Energy_Bin_145 <= s_Energy_Bin_145;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_145 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_145;  
 
  
  Energy_Bin_146 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_146   <=  (others =>'0');
		Energy_Bin_Rdy_146 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E146_C1_L and PEAK_C1 <= s_E146_C1_H and Bin_OR = '0') then
         s_Energy_Bin_146 <= s_Energy_Bin_146 +'1';
		 Energy_Bin_Rdy_146 <= '1';
		else
		 s_Energy_Bin_146 <= s_Energy_Bin_146;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_146 <= '0';
      end if;
    end if;
  end process  Energy_Bin_146;   
  
 Energy_Bin_147 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_147   <=  (others =>'0');
		Energy_Bin_Rdy_147 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E147_C1_L and PEAK_C1 <= s_E147_C1_H and Bin_OR = '0') then
         s_Energy_Bin_147 <= s_Energy_Bin_147 +'1';
		 Energy_Bin_Rdy_147 <= '1';
		else
		 s_Energy_Bin_147 <= s_Energy_Bin_147;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_147 <= '0';
      end if;
    end if;
  end process  Energy_Bin_147;   
  
  Energy_Bin_148 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_148   <=  (others =>'0');
		Energy_Bin_Rdy_148 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E148_C1_L and PEAK_C1 <= s_E148_C1_H and Bin_OR = '0') then
         s_Energy_Bin_148 <= s_Energy_Bin_148 +'1';
		 Energy_Bin_Rdy_148 <= '1';
		else
		 s_Energy_Bin_148 <= s_Energy_Bin_148;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_148 <= '0';
      end if;
    end if;
  end process  Energy_Bin_148;   
  
  Energy_Bin_149 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_149   <=  (others =>'0');
		Energy_Bin_Rdy_149 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E149_C1_L and PEAK_C1 <= s_E149_C1_H and Bin_OR = '0') then
         s_Energy_Bin_149 <= s_Energy_Bin_149 +'1';
		 Energy_Bin_Rdy_149 <= '1';
		else
		 s_Energy_Bin_149 <= s_Energy_Bin_149;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_149 <= '0';
      end if;
    end if;
  end process  Energy_Bin_149;          
  
  
     Energy_Bin_150 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_150   <=  (others =>'0');
		Energy_Bin_Rdy_150 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E150_C1_L and PEAK_C1 <= s_E150_C1_H and Bin_OR = '0') then
         s_Energy_Bin_150 <= s_Energy_Bin_150 +'1';
		 Energy_Bin_Rdy_150 <= '1';
		else
		 s_Energy_Bin_150 <= s_Energy_Bin_150;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_150 <= '0';
      end if;
    end if;
  end process  Energy_Bin_150;    
  
  Energy_Bin_151 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_151   <=  (others =>'0');
		Energy_Bin_Rdy_151 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E151_C1_L and PEAK_C1 <= s_E151_C1_H and Bin_OR = '0') then
         s_Energy_Bin_151 <= s_Energy_Bin_151 +'1';
		 Energy_Bin_Rdy_151 <= '1';
		else
		 s_Energy_Bin_151 <= s_Energy_Bin_151;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_151 <= '0';
      end if;
    end if;
  end process  Energy_Bin_151;   
  
  Energy_Bin_152 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_152   <=  (others =>'0');
	    Energy_Bin_Rdy_152 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E152_C1_L and PEAK_C1 <= s_E152_C1_H and Bin_OR = '0') then
         s_Energy_Bin_152 <= s_Energy_Bin_152 +'1';
		 Energy_Bin_Rdy_152 <= '1';
		else
		 s_Energy_Bin_152 <= s_Energy_Bin_152;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_152 <= '0';
      end if;
    end if;
  end process  Energy_Bin_152;   
  
  Energy_Bin_153 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_153   <=  (others =>'0');
	    Energy_Bin_Rdy_153 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E153_C1_L and PEAK_C1 <= s_E153_C1_H and Bin_OR = '0') then
         s_Energy_Bin_153 <= s_Energy_Bin_153 +'1';
		 Energy_Bin_Rdy_153 <= '1';
		else
		 s_Energy_Bin_153 <= s_Energy_Bin_153;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_153 <= '0';
      end if;
    end if;
  end process  Energy_Bin_153;   
  
  Energy_Bin_154 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_154   <=  (others =>'0');
		Energy_Bin_Rdy_154 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E154_C1_L and PEAK_C1 <= s_E154_C1_H and Bin_OR = '0') then
         s_Energy_Bin_154 <= s_Energy_Bin_154 +'1';
		 Energy_Bin_Rdy_154 <= '1';
		else
		 s_Energy_Bin_154 <= s_Energy_Bin_154;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_154 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_154;   
 
 
  Energy_Bin_155 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_155   <=  (others =>'0');
		Energy_Bin_Rdy_155 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E155_C1_L and PEAK_C1 <= s_E155_C1_H and Bin_OR = '0') then
         s_Energy_Bin_155 <= s_Energy_Bin_155 +'1';
		 Energy_Bin_Rdy_155 <= '1';
		else
		 s_Energy_Bin_155 <= s_Energy_Bin_155;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_155 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_155;  
 
  
  Energy_Bin_156 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_156   <=  (others =>'0');
		Energy_Bin_Rdy_156 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E156_C1_L and PEAK_C1 <= s_E156_C1_H and Bin_OR = '0') then
         s_Energy_Bin_156 <= s_Energy_Bin_156 +'1';
		 Energy_Bin_Rdy_156 <= '1';
		else
		 s_Energy_Bin_156 <= s_Energy_Bin_156;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_156 <= '0';
      end if;
    end if;
  end process  Energy_Bin_156;   
  
 Energy_Bin_157 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_157   <=  (others =>'0');
		Energy_Bin_Rdy_157 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E157_C1_L and PEAK_C1 <= s_E157_C1_H and Bin_OR = '0') then
         s_Energy_Bin_157 <= s_Energy_Bin_157 +'1';
		 Energy_Bin_Rdy_157 <= '1';
		else
		 s_Energy_Bin_157 <= s_Energy_Bin_157;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_157 <= '0';
      end if;
    end if;
  end process  Energy_Bin_157;   
  
  Energy_Bin_158 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_158   <=  (others =>'0');
		Energy_Bin_Rdy_158 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E158_C1_L and PEAK_C1 <= s_E158_C1_H and Bin_OR = '0') then
         s_Energy_Bin_158 <= s_Energy_Bin_158 +'1';
		 Energy_Bin_Rdy_158 <= '1';
		else
		 s_Energy_Bin_158 <= s_Energy_Bin_158;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_158 <= '0';
      end if;
    end if;
  end process  Energy_Bin_158;   
  
  Energy_Bin_159 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_159   <=  (others =>'0');
		Energy_Bin_Rdy_159 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E159_C1_L and PEAK_C1 <= s_E159_C1_H and Bin_OR = '0') then
         s_Energy_Bin_159 <= s_Energy_Bin_159 +'1';
		 Energy_Bin_Rdy_159 <= '1';
		else
		 s_Energy_Bin_159 <= s_Energy_Bin_159;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_159 <= '0';
      end if;
    end if;
  end process  Energy_Bin_159;           
  
     Energy_Bin_160 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_160   <=  (others =>'0');
		Energy_Bin_Rdy_160 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E160_C1_L and PEAK_C1 <= s_E160_C1_H and Bin_OR = '0') then
         s_Energy_Bin_160 <= s_Energy_Bin_160 +'1';
		 Energy_Bin_Rdy_160 <= '1';
		else
		 s_Energy_Bin_160 <= s_Energy_Bin_160;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_160 <= '0';
      end if;
    end if;
  end process  Energy_Bin_160;    
  
  Energy_Bin_161 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_161   <=  (others =>'0');
		Energy_Bin_Rdy_161 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E161_C1_L and PEAK_C1 <= s_E161_C1_H and Bin_OR = '0') then
         s_Energy_Bin_161 <= s_Energy_Bin_161 +'1';
		 Energy_Bin_Rdy_161 <= '1';
		else
		 s_Energy_Bin_161 <= s_Energy_Bin_161;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_161 <= '0';
      end if;
    end if;
  end process  Energy_Bin_161;   
  
  Energy_Bin_162 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_162   <=  (others =>'0');
	    Energy_Bin_Rdy_162 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E162_C1_L and PEAK_C1 <= s_E162_C1_H and Bin_OR = '0') then
         s_Energy_Bin_162 <= s_Energy_Bin_162 +'1';
		 Energy_Bin_Rdy_162 <= '1';
		else
		 s_Energy_Bin_162 <= s_Energy_Bin_162;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_162 <= '0';
      end if;
    end if;
  end process  Energy_Bin_162;   
  
  Energy_Bin_163 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_163   <=  (others =>'0');
	    Energy_Bin_Rdy_163 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E163_C1_L and PEAK_C1 <= s_E163_C1_H and Bin_OR = '0') then
         s_Energy_Bin_163 <= s_Energy_Bin_163 +'1';
		 Energy_Bin_Rdy_163 <= '1';
		else
		 s_Energy_Bin_163 <= s_Energy_Bin_163;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_163 <= '0';
      end if;
    end if;
  end process  Energy_Bin_163;   
  
  Energy_Bin_164 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_164   <=  (others =>'0');
		Energy_Bin_Rdy_164 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E164_C1_L and PEAK_C1 <= s_E164_C1_H and Bin_OR = '0') then
         s_Energy_Bin_164 <= s_Energy_Bin_164 +'1';
		 Energy_Bin_Rdy_164 <= '1';
		else
		 s_Energy_Bin_164 <= s_Energy_Bin_164;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_164 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_164;   
 
 
  Energy_Bin_165 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_165   <=  (others =>'0');
		Energy_Bin_Rdy_165 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E165_C1_L and PEAK_C1 <= s_E165_C1_H and Bin_OR = '0') then
         s_Energy_Bin_165 <= s_Energy_Bin_165 +'1';
		 Energy_Bin_Rdy_165 <= '1';
		else
		 s_Energy_Bin_165 <= s_Energy_Bin_165;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_165 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_165;  
 
  
  Energy_Bin_166 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_166   <=  (others =>'0');
		Energy_Bin_Rdy_166 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E166_C1_L and PEAK_C1 <= s_E166_C1_H and Bin_OR = '0') then
         s_Energy_Bin_166 <= s_Energy_Bin_166 +'1';
		 Energy_Bin_Rdy_166 <= '1';
		else
		 s_Energy_Bin_166 <= s_Energy_Bin_166;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_166 <= '0';
      end if;
    end if;
  end process  Energy_Bin_166;   
  
 Energy_Bin_167 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_167   <=  (others =>'0');
		Energy_Bin_Rdy_167 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E167_C1_L and PEAK_C1 <= s_E167_C1_H and Bin_OR = '0') then
         s_Energy_Bin_167 <= s_Energy_Bin_167 +'1';
		 Energy_Bin_Rdy_167 <= '1';
		else
		 s_Energy_Bin_167 <= s_Energy_Bin_167;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_167 <= '0';
      end if;
    end if;
  end process  Energy_Bin_167;   
  
  Energy_Bin_168 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_168   <=  (others =>'0');
		Energy_Bin_Rdy_168 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E168_C1_L and PEAK_C1 <= s_E168_C1_H and Bin_OR = '0') then
         s_Energy_Bin_168 <= s_Energy_Bin_168 +'1';
		 Energy_Bin_Rdy_168 <= '1';
		else
		 s_Energy_Bin_168 <= s_Energy_Bin_168;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_168 <= '0';
      end if;
    end if;
  end process  Energy_Bin_168;   
  
  Energy_Bin_169 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_169   <=  (others =>'0');
		Energy_Bin_Rdy_169 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E169_C1_L and PEAK_C1 <= s_E169_C1_H and Bin_OR = '0') then
         s_Energy_Bin_169 <= s_Energy_Bin_169 +'1';
		 Energy_Bin_Rdy_169 <= '1';
		else
		 s_Energy_Bin_169 <= s_Energy_Bin_169;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_169 <= '0';
      end if;
    end if;
  end process  Energy_Bin_169;         
  
     Energy_Bin_170 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_170   <=  (others =>'0');
		Energy_Bin_Rdy_170 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E170_C1_L and PEAK_C1 <= s_E170_C1_H and Bin_OR = '0') then
         s_Energy_Bin_170 <= s_Energy_Bin_170 +'1';
		 Energy_Bin_Rdy_170 <= '1';
		else
		 s_Energy_Bin_170 <= s_Energy_Bin_170;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_170 <= '0';
      end if;
    end if;
  end process  Energy_Bin_170;    
  
  Energy_Bin_171 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_171   <=  (others =>'0');
		Energy_Bin_Rdy_171 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E171_C1_L and PEAK_C1 <= s_E171_C1_H and Bin_OR = '0') then
         s_Energy_Bin_171 <= s_Energy_Bin_171 +'1';
		 Energy_Bin_Rdy_171 <= '1';
		else
		 s_Energy_Bin_171 <= s_Energy_Bin_171;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_171 <= '0';
      end if;
    end if;
  end process  Energy_Bin_171;   
  
  Energy_Bin_172 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_172   <=  (others =>'0');
	    Energy_Bin_Rdy_172 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E172_C1_L and PEAK_C1 <= s_E172_C1_H and Bin_OR = '0') then
         s_Energy_Bin_172 <= s_Energy_Bin_172 +'1';
		 Energy_Bin_Rdy_172 <= '1';
		else
		 s_Energy_Bin_172 <= s_Energy_Bin_172;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_172 <= '0';
      end if;
    end if;
  end process  Energy_Bin_172;   
  
  Energy_Bin_173 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_173   <=  (others =>'0');
	    Energy_Bin_Rdy_173 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E173_C1_L and PEAK_C1 <= s_E173_C1_H and Bin_OR = '0') then
         s_Energy_Bin_173 <= s_Energy_Bin_173 +'1';
		 Energy_Bin_Rdy_173 <= '1';
		else
		 s_Energy_Bin_173 <= s_Energy_Bin_173;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_173 <= '0';
      end if;
    end if;
  end process  Energy_Bin_173;   
  
  Energy_Bin_174 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_174   <=  (others =>'0');
		Energy_Bin_Rdy_174 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E174_C1_L and PEAK_C1 <= s_E174_C1_H and Bin_OR = '0') then
         s_Energy_Bin_174 <= s_Energy_Bin_174 +'1';
		 Energy_Bin_Rdy_174 <= '1';
		else
		 s_Energy_Bin_174 <= s_Energy_Bin_174;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_174 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_174;   
 
 
  Energy_Bin_175 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_175   <=  (others =>'0');
		Energy_Bin_Rdy_175 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E175_C1_L and PEAK_C1 <= s_E175_C1_H and Bin_OR = '0') then
         s_Energy_Bin_175 <= s_Energy_Bin_175 +'1';
		 Energy_Bin_Rdy_175 <= '1';
		else
		 s_Energy_Bin_175 <= s_Energy_Bin_175;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_175 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_175;  
 
  
  Energy_Bin_176 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_176   <=  (others =>'0');
		Energy_Bin_Rdy_176 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E176_C1_L and PEAK_C1 <= s_E176_C1_H and Bin_OR = '0') then
         s_Energy_Bin_176 <= s_Energy_Bin_176 +'1';
		 Energy_Bin_Rdy_176 <= '1';
		else
		 s_Energy_Bin_176 <= s_Energy_Bin_176;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_176 <= '0';
      end if;
    end if;
  end process  Energy_Bin_176;   
  
 Energy_Bin_177 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_177   <=  (others =>'0');
		Energy_Bin_Rdy_177 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E177_C1_L and PEAK_C1 <= s_E177_C1_H and Bin_OR = '0') then
         s_Energy_Bin_177 <= s_Energy_Bin_177 +'1';
		 Energy_Bin_Rdy_177 <= '1';
		else
		 s_Energy_Bin_177 <= s_Energy_Bin_177;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_177 <= '0';
      end if;
    end if;
  end process  Energy_Bin_177;   
  
  Energy_Bin_178 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_178   <=  (others =>'0');
		Energy_Bin_Rdy_178 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E178_C1_L and PEAK_C1 <= s_E178_C1_H and Bin_OR = '0') then
         s_Energy_Bin_178 <= s_Energy_Bin_178 +'1';
		 Energy_Bin_Rdy_178 <= '1';
		else
		 s_Energy_Bin_178 <= s_Energy_Bin_178;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_178 <= '0';
      end if;
    end if;
  end process  Energy_Bin_178;   
  
  Energy_Bin_179 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_179   <=  (others =>'0');
		Energy_Bin_Rdy_179 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E179_C1_L and PEAK_C1 <= s_E179_C1_H and Bin_OR = '0') then
         s_Energy_Bin_179 <= s_Energy_Bin_179 +'1';
		 Energy_Bin_Rdy_179 <= '1';
		else
		 s_Energy_Bin_179 <= s_Energy_Bin_179;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_179 <= '0';
      end if;
    end if;
  end process  Energy_Bin_179;       
  
     Energy_Bin_180 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_180   <=  (others =>'0');
		Energy_Bin_Rdy_180 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E180_C1_L and PEAK_C1 <= s_E180_C1_H and Bin_OR = '0') then
         s_Energy_Bin_180 <= s_Energy_Bin_180 +'1';
		 Energy_Bin_Rdy_180 <= '1';
		else
		 s_Energy_Bin_180 <= s_Energy_Bin_180;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_180 <= '0';
      end if;
    end if;
  end process  Energy_Bin_180;    
  
  Energy_Bin_181 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_181   <=  (others =>'0');
		Energy_Bin_Rdy_181 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E181_C1_L and PEAK_C1 <= s_E181_C1_H and Bin_OR = '0') then
         s_Energy_Bin_181 <= s_Energy_Bin_181 +'1';
		 Energy_Bin_Rdy_181 <= '1';
		else
		 s_Energy_Bin_181 <= s_Energy_Bin_181;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_181 <= '0';
      end if;
    end if;
  end process  Energy_Bin_181;   
  
  Energy_Bin_182 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_182   <=  (others =>'0');
	    Energy_Bin_Rdy_182 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E182_C1_L and PEAK_C1 <= s_E182_C1_H and Bin_OR = '0') then
         s_Energy_Bin_182 <= s_Energy_Bin_182 +'1';
		 Energy_Bin_Rdy_182 <= '1';
		else
		 s_Energy_Bin_182 <= s_Energy_Bin_182;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_182 <= '0';
      end if;
    end if;
  end process  Energy_Bin_182;   
  
  Energy_Bin_183 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_183   <=  (others =>'0');
	    Energy_Bin_Rdy_183 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E183_C1_L and PEAK_C1 <= s_E183_C1_H and Bin_OR = '0') then
         s_Energy_Bin_183 <= s_Energy_Bin_183 +'1';
		 Energy_Bin_Rdy_183 <= '1';
		else
		 s_Energy_Bin_183 <= s_Energy_Bin_183;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_183 <= '0';
      end if;
    end if;
  end process  Energy_Bin_183;   
  
  Energy_Bin_184 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_184   <=  (others =>'0');
		Energy_Bin_Rdy_184 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E184_C1_L and PEAK_C1 <= s_E184_C1_H and Bin_OR = '0') then
         s_Energy_Bin_184 <= s_Energy_Bin_184 +'1';
		 Energy_Bin_Rdy_184 <= '1';
		else
		 s_Energy_Bin_184 <= s_Energy_Bin_184;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_184 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_184;   
 
 
  Energy_Bin_185 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_185   <=  (others =>'0');
		Energy_Bin_Rdy_185 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E185_C1_L and PEAK_C1 <= s_E185_C1_H and Bin_OR = '0') then
         s_Energy_Bin_185 <= s_Energy_Bin_185 +'1';
		 Energy_Bin_Rdy_185 <= '1';
		else
		 s_Energy_Bin_185 <= s_Energy_Bin_185;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_185 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_185;  
 
  
  Energy_Bin_186 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_186   <=  (others =>'0');
		Energy_Bin_Rdy_186 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E186_C1_L and PEAK_C1 <= s_E186_C1_H and Bin_OR = '0') then
         s_Energy_Bin_186 <= s_Energy_Bin_186 +'1';
		 Energy_Bin_Rdy_186 <= '1';
		else
		 s_Energy_Bin_186 <= s_Energy_Bin_186;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_186 <= '0';
      end if;
    end if;
  end process  Energy_Bin_186;   
  
 Energy_Bin_187 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_187   <=  (others =>'0');
		Energy_Bin_Rdy_187 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E187_C1_L and PEAK_C1 <= s_E187_C1_H and Bin_OR = '0') then
         s_Energy_Bin_187 <= s_Energy_Bin_187 +'1';
		 Energy_Bin_Rdy_187 <= '1';
		else
		 s_Energy_Bin_187 <= s_Energy_Bin_187;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_187 <= '0';
      end if;
    end if;
  end process  Energy_Bin_187;   
  
  Energy_Bin_188 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_188   <=  (others =>'0');
		Energy_Bin_Rdy_188 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E188_C1_L and PEAK_C1 <= s_E188_C1_H and Bin_OR = '0') then
         s_Energy_Bin_188 <= s_Energy_Bin_188 +'1';
		 Energy_Bin_Rdy_188 <= '1';
		else
		 s_Energy_Bin_188 <= s_Energy_Bin_188;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_188 <= '0';
      end if;
    end if;
  end process  Energy_Bin_188;   
  
  Energy_Bin_189 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_189   <=  (others =>'0');
		Energy_Bin_Rdy_189 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E189_C1_L and PEAK_C1 <= s_E189_C1_H and Bin_OR = '0') then
         s_Energy_Bin_189 <= s_Energy_Bin_189 +'1';
		 Energy_Bin_Rdy_189 <= '1';
		else
		 s_Energy_Bin_189 <= s_Energy_Bin_189;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_189 <= '0';
      end if;
    end if;
  end process  Energy_Bin_189;      
  
     Energy_Bin_190 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_190   <=  (others =>'0');
		Energy_Bin_Rdy_190 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E190_C1_L and PEAK_C1 <= s_E190_C1_H and Bin_OR = '0') then
         s_Energy_Bin_190 <= s_Energy_Bin_190 +'1';
		 Energy_Bin_Rdy_190 <= '1';
		else
		 s_Energy_Bin_190 <= s_Energy_Bin_190;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_190 <= '0';
      end if;
    end if;
  end process  Energy_Bin_190;    
  
  Energy_Bin_191 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_191   <=  (others =>'0');
		Energy_Bin_Rdy_191 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E191_C1_L and PEAK_C1 <= s_E191_C1_H and Bin_OR = '0') then
         s_Energy_Bin_191 <= s_Energy_Bin_191 +'1';
		 Energy_Bin_Rdy_191 <= '1';
		else
		 s_Energy_Bin_191 <= s_Energy_Bin_191;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_191 <= '0';
      end if;
    end if;
  end process  Energy_Bin_191;   
  
  Energy_Bin_192 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_192   <=  (others =>'0');
	    Energy_Bin_Rdy_192 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E192_C1_L and PEAK_C1 <= s_E192_C1_H and Bin_OR = '0') then
         s_Energy_Bin_192 <= s_Energy_Bin_192 +'1';
		 Energy_Bin_Rdy_192 <= '1';
		else
		 s_Energy_Bin_192 <= s_Energy_Bin_192;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_192 <= '0';
      end if;
    end if;
  end process  Energy_Bin_192;   
  
  Energy_Bin_193 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_193   <=  (others =>'0');
	    Energy_Bin_Rdy_193 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E193_C1_L and PEAK_C1 <= s_E193_C1_H and Bin_OR = '0') then
         s_Energy_Bin_193 <= s_Energy_Bin_193 +'1';
		 Energy_Bin_Rdy_193 <= '1';
		else
		 s_Energy_Bin_193 <= s_Energy_Bin_193;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_193 <= '0';
      end if;
    end if;
  end process  Energy_Bin_193;   
  
  Energy_Bin_194 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_194   <=  (others =>'0');
		Energy_Bin_Rdy_194 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E194_C1_L and PEAK_C1 <= s_E194_C1_H and Bin_OR = '0') then
         s_Energy_Bin_194 <= s_Energy_Bin_194 +'1';
		 Energy_Bin_Rdy_194 <= '1';
		else
		 s_Energy_Bin_194 <= s_Energy_Bin_194;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_194 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_194;   
 
 
  Energy_Bin_195 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_195   <=  (others =>'0');
		Energy_Bin_Rdy_195 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E195_C1_L and PEAK_C1 <= s_E195_C1_H and Bin_OR = '0') then
         s_Energy_Bin_195 <= s_Energy_Bin_195 +'1';
		 Energy_Bin_Rdy_195 <= '1';
		else
		 s_Energy_Bin_195 <= s_Energy_Bin_195;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_195 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_195;  
 
  
  Energy_Bin_196 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_196   <=  (others =>'0');
		Energy_Bin_Rdy_196 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E196_C1_L and PEAK_C1 <= s_E196_C1_H and Bin_OR = '0') then
         s_Energy_Bin_196 <= s_Energy_Bin_196 +'1';
		 Energy_Bin_Rdy_196 <= '1';
		else
		 s_Energy_Bin_196 <= s_Energy_Bin_196;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_196 <= '0';
      end if;
    end if;
  end process  Energy_Bin_196;   
  
 Energy_Bin_197 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_197   <=  (others =>'0');
		Energy_Bin_Rdy_197 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E197_C1_L and PEAK_C1 <= s_E197_C1_H and Bin_OR = '0') then
         s_Energy_Bin_197 <= s_Energy_Bin_197 +'1';
		 Energy_Bin_Rdy_197 <= '1';
		else
		 s_Energy_Bin_197 <= s_Energy_Bin_197;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_197 <= '0';
      end if;
    end if;
  end process  Energy_Bin_197;   
  
  Energy_Bin_198 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_198   <=  (others =>'0');
		Energy_Bin_Rdy_198 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E198_C1_L and PEAK_C1 <= s_E198_C1_H and Bin_OR = '0') then
         s_Energy_Bin_198 <= s_Energy_Bin_198 +'1';
		 Energy_Bin_Rdy_198 <= '1';
		else
		 s_Energy_Bin_198 <= s_Energy_Bin_198;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_198 <= '0';
      end if;
    end if;
  end process  Energy_Bin_198;   
  
  Energy_Bin_199 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_199   <=  (others =>'0');
		Energy_Bin_Rdy_199 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E199_C1_L and PEAK_C1 <= s_E199_C1_H and Bin_OR = '0') then
         s_Energy_Bin_199 <= s_Energy_Bin_199 +'1';
		 Energy_Bin_Rdy_199 <= '1';
		else
		 s_Energy_Bin_199 <= s_Energy_Bin_199;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_199 <= '0';
      end if;
    end if;
  end process  Energy_Bin_199;      
    
     Energy_Bin_200 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_200   <=  (others =>'0');
		Energy_Bin_Rdy_200 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E200_C1_L and PEAK_C1 <= s_E200_C1_H and Bin_OR = '0') then
         s_Energy_Bin_200 <= s_Energy_Bin_200 +'1';
		 Energy_Bin_Rdy_200 <= '1';
		else
		 s_Energy_Bin_200 <= s_Energy_Bin_200;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_200 <= '0';
      end if;
    end if;
  end process  Energy_Bin_200;    
  
  Energy_Bin_201 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_201   <=  (others =>'0');
		Energy_Bin_Rdy_201 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E201_C1_L and PEAK_C1 <= s_E201_C1_H and Bin_OR = '0') then
         s_Energy_Bin_201 <= s_Energy_Bin_201 +'1';
		 Energy_Bin_Rdy_201 <= '1';
		else
		 s_Energy_Bin_201 <= s_Energy_Bin_201;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_201 <= '0';
      end if;
    end if;
  end process  Energy_Bin_201;   
  
  Energy_Bin_202 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_202   <=  (others =>'0');
	    Energy_Bin_Rdy_202 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E202_C1_L and PEAK_C1 <= s_E202_C1_H and Bin_OR = '0') then
         s_Energy_Bin_202 <= s_Energy_Bin_202 +'1';
		 Energy_Bin_Rdy_202 <= '1';
		else
		 s_Energy_Bin_202 <= s_Energy_Bin_202;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_202 <= '0';
      end if;
    end if;
  end process  Energy_Bin_202;   
  
  Energy_Bin_203 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_203   <=  (others =>'0');
	    Energy_Bin_Rdy_203 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E203_C1_L and PEAK_C1 <= s_E203_C1_H and Bin_OR = '0') then
         s_Energy_Bin_203 <= s_Energy_Bin_203 +'1';
		 Energy_Bin_Rdy_203 <= '1';
		else
		 s_Energy_Bin_203 <= s_Energy_Bin_203;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_203 <= '0';
      end if;
    end if;
  end process  Energy_Bin_203;   
  
  Energy_Bin_204 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_204   <=  (others =>'0');
		Energy_Bin_Rdy_204 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E204_C1_L and PEAK_C1 <= s_E204_C1_H and Bin_OR = '0') then
         s_Energy_Bin_204 <= s_Energy_Bin_204 +'1';
		 Energy_Bin_Rdy_204 <= '1';
		else
		 s_Energy_Bin_204 <= s_Energy_Bin_204;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_204 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_204;   
 
 
  Energy_Bin_205 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_205   <=  (others =>'0');
		Energy_Bin_Rdy_205 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E205_C1_L and PEAK_C1 <= s_E205_C1_H and Bin_OR = '0') then
         s_Energy_Bin_205 <= s_Energy_Bin_205 +'1';
		 Energy_Bin_Rdy_205 <= '1';
		else
		 s_Energy_Bin_205 <= s_Energy_Bin_205;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_205 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_205;  
 
  
  Energy_Bin_206 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_206   <=  (others =>'0');
		Energy_Bin_Rdy_206 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E206_C1_L and PEAK_C1 <= s_E206_C1_H and Bin_OR = '0') then
         s_Energy_Bin_206 <= s_Energy_Bin_206 +'1';
		 Energy_Bin_Rdy_206 <= '1';
		else
		 s_Energy_Bin_206 <= s_Energy_Bin_206;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_206 <= '0';
      end if;
    end if;
  end process  Energy_Bin_206;   
  
 Energy_Bin_207 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_207   <=  (others =>'0');
		Energy_Bin_Rdy_207 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E207_C1_L and PEAK_C1 <= s_E207_C1_H and Bin_OR = '0') then
         s_Energy_Bin_207 <= s_Energy_Bin_207 +'1';
		 Energy_Bin_Rdy_207 <= '1';
		else
		 s_Energy_Bin_207 <= s_Energy_Bin_207;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_207 <= '0';
      end if;
    end if;
  end process  Energy_Bin_207;   
  
  Energy_Bin_208 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_208   <=  (others =>'0');
		Energy_Bin_Rdy_208 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E208_C1_L and PEAK_C1 <= s_E208_C1_H and Bin_OR = '0') then
         s_Energy_Bin_208 <= s_Energy_Bin_208 +'1';
		 Energy_Bin_Rdy_208 <= '1';
		else
		 s_Energy_Bin_208 <= s_Energy_Bin_208;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_208 <= '0';
      end if;
    end if;
  end process  Energy_Bin_208;   
  
  Energy_Bin_209 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_209   <=  (others =>'0');
		Energy_Bin_Rdy_209 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E209_C1_L and PEAK_C1 <= s_E209_C1_H and Bin_OR = '0') then
         s_Energy_Bin_209 <= s_Energy_Bin_209 +'1';
		 Energy_Bin_Rdy_209 <= '1';
		else
		 s_Energy_Bin_209 <= s_Energy_Bin_209;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_209 <= '0';
      end if;
    end if;
  end process  Energy_Bin_209;      
  
     Energy_Bin_210 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_210   <=  (others =>'0');
		Energy_Bin_Rdy_210 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E210_C1_L and PEAK_C1 <= s_E210_C1_H and Bin_OR = '0') then
         s_Energy_Bin_210 <= s_Energy_Bin_210 +'1';
		 Energy_Bin_Rdy_210 <= '1';
		else
		 s_Energy_Bin_210 <= s_Energy_Bin_210;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_210 <= '0';
      end if;
    end if;
  end process  Energy_Bin_210;    
  
  Energy_Bin_211 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_211   <=  (others =>'0');
		Energy_Bin_Rdy_211 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E211_C1_L and PEAK_C1 <= s_E211_C1_H and Bin_OR = '0') then
         s_Energy_Bin_211 <= s_Energy_Bin_211 +'1';
		 Energy_Bin_Rdy_211 <= '1';
		else
		 s_Energy_Bin_211 <= s_Energy_Bin_211;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_211 <= '0';
      end if;
    end if;
  end process  Energy_Bin_211;   
  
  Energy_Bin_212 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_212   <=  (others =>'0');
	    Energy_Bin_Rdy_212 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E212_C1_L and PEAK_C1 <= s_E212_C1_H and Bin_OR = '0') then
         s_Energy_Bin_212 <= s_Energy_Bin_212 +'1';
		 Energy_Bin_Rdy_212 <= '1';
		else
		 s_Energy_Bin_212 <= s_Energy_Bin_212;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_212 <= '0';
      end if;
    end if;
  end process  Energy_Bin_212;   
  
  Energy_Bin_213 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_213   <=  (others =>'0');
	    Energy_Bin_Rdy_213 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E213_C1_L and PEAK_C1 <= s_E213_C1_H and Bin_OR = '0') then
         s_Energy_Bin_213 <= s_Energy_Bin_213 +'1';
		 Energy_Bin_Rdy_213 <= '1';
		else
		 s_Energy_Bin_213 <= s_Energy_Bin_213;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_213 <= '0';
      end if;
    end if;
  end process  Energy_Bin_213;   
  
  Energy_Bin_214 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_214   <=  (others =>'0');
		Energy_Bin_Rdy_214 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E214_C1_L and PEAK_C1 <= s_E214_C1_H and Bin_OR = '0') then
         s_Energy_Bin_214 <= s_Energy_Bin_214 +'1';
		 Energy_Bin_Rdy_214 <= '1';
		else
		 s_Energy_Bin_214 <= s_Energy_Bin_214;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_214 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_214;   
 
 
  Energy_Bin_215 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_215   <=  (others =>'0');
		Energy_Bin_Rdy_215 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E215_C1_L and PEAK_C1 <= s_E215_C1_H and Bin_OR = '0') then
         s_Energy_Bin_215 <= s_Energy_Bin_215 +'1';
		 Energy_Bin_Rdy_215 <= '1';
		else
		 s_Energy_Bin_215 <= s_Energy_Bin_215;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_215 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_215;  
 
  
  Energy_Bin_216 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_216   <=  (others =>'0');
		Energy_Bin_Rdy_216 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E216_C1_L and PEAK_C1 <= s_E216_C1_H and Bin_OR = '0') then
         s_Energy_Bin_216 <= s_Energy_Bin_216 +'1';
		 Energy_Bin_Rdy_216 <= '1';
		else
		 s_Energy_Bin_216 <= s_Energy_Bin_216;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_216 <= '0';
      end if;
    end if;
  end process  Energy_Bin_216;   
  
 Energy_Bin_217 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_217   <=  (others =>'0');
		Energy_Bin_Rdy_217 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E217_C1_L and PEAK_C1 <= s_E217_C1_H and Bin_OR = '0') then
         s_Energy_Bin_217 <= s_Energy_Bin_217 +'1';
		 Energy_Bin_Rdy_217 <= '1';
		else
		 s_Energy_Bin_217 <= s_Energy_Bin_217;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_217 <= '0';
      end if;
    end if;
  end process  Energy_Bin_217;   
  
  Energy_Bin_218 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_218   <=  (others =>'0');
		Energy_Bin_Rdy_218 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E218_C1_L and PEAK_C1 <= s_E218_C1_H and Bin_OR = '0') then
         s_Energy_Bin_218 <= s_Energy_Bin_218 +'1';
		 Energy_Bin_Rdy_218 <= '1';
		else
		 s_Energy_Bin_218 <= s_Energy_Bin_218;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_218 <= '0';
      end if;
    end if;
  end process  Energy_Bin_218;   
  
  Energy_Bin_219 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_219   <=  (others =>'0');
		Energy_Bin_Rdy_219 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E219_C1_L and PEAK_C1 <= s_E219_C1_H and Bin_OR = '0') then
         s_Energy_Bin_219 <= s_Energy_Bin_219 +'1';
		 Energy_Bin_Rdy_219 <= '1';
		else
		 s_Energy_Bin_219 <= s_Energy_Bin_219;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_219 <= '0';
      end if;
    end if;
  end process  Energy_Bin_219;       
  
     Energy_Bin_220 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_220   <=  (others =>'0');
		Energy_Bin_Rdy_220 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E220_C1_L and PEAK_C1 <= s_E220_C1_H and Bin_OR = '0') then
         s_Energy_Bin_220 <= s_Energy_Bin_220 +'1';
		 Energy_Bin_Rdy_220 <= '1';
		else
		 s_Energy_Bin_220 <= s_Energy_Bin_220;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_220 <= '0';
      end if;
    end if;
  end process  Energy_Bin_220;    
  
  Energy_Bin_221 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_221   <=  (others =>'0');
		Energy_Bin_Rdy_221 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E221_C1_L and PEAK_C1 <= s_E221_C1_H and Bin_OR = '0') then
         s_Energy_Bin_221 <= s_Energy_Bin_221 +'1';
		 Energy_Bin_Rdy_221 <= '1';
		else
		 s_Energy_Bin_221 <= s_Energy_Bin_221;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_221 <= '0';
      end if;
    end if;
  end process  Energy_Bin_221;   
  
  Energy_Bin_222 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_222   <=  (others =>'0');
	    Energy_Bin_Rdy_222 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E222_C1_L and PEAK_C1 <= s_E222_C1_H and Bin_OR = '0') then
         s_Energy_Bin_222 <= s_Energy_Bin_222 +'1';
		 Energy_Bin_Rdy_222 <= '1';
		else
		 s_Energy_Bin_222 <= s_Energy_Bin_222;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_222 <= '0';
      end if;
    end if;
  end process  Energy_Bin_222;   
  
  Energy_Bin_223 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_223   <=  (others =>'0');
	    Energy_Bin_Rdy_223 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E223_C1_L and PEAK_C1 <= s_E223_C1_H and Bin_OR = '0') then
         s_Energy_Bin_223 <= s_Energy_Bin_223 +'1';
		 Energy_Bin_Rdy_223 <= '1';
		else
		 s_Energy_Bin_223 <= s_Energy_Bin_223;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_223 <= '0';
      end if;
    end if;
  end process  Energy_Bin_223;   
  
  Energy_Bin_224 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_224   <=  (others =>'0');
		Energy_Bin_Rdy_224 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E224_C1_L and PEAK_C1 <= s_E224_C1_H and Bin_OR = '0') then
         s_Energy_Bin_224 <= s_Energy_Bin_224 +'1';
		 Energy_Bin_Rdy_224 <= '1';
		else
		 s_Energy_Bin_224 <= s_Energy_Bin_224;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_224 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_224;   
 
 
  Energy_Bin_225 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_225   <=  (others =>'0');
		Energy_Bin_Rdy_225 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E225_C1_L and PEAK_C1 <= s_E225_C1_H and Bin_OR = '0') then
         s_Energy_Bin_225 <= s_Energy_Bin_225 +'1';
		 Energy_Bin_Rdy_225 <= '1';
		else
		 s_Energy_Bin_225 <= s_Energy_Bin_225;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_225 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_225;  
 
  
  Energy_Bin_226 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_226   <=  (others =>'0');
		Energy_Bin_Rdy_226 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E226_C1_L and PEAK_C1 <= s_E226_C1_H and Bin_OR = '0') then
         s_Energy_Bin_226 <= s_Energy_Bin_226 +'1';
		 Energy_Bin_Rdy_226 <= '1';
		else
		 s_Energy_Bin_226 <= s_Energy_Bin_226;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_226 <= '0';
      end if;
    end if;
  end process  Energy_Bin_226;   
  
 Energy_Bin_227 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_227   <=  (others =>'0');
		Energy_Bin_Rdy_227 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E227_C1_L and PEAK_C1 <= s_E227_C1_H and Bin_OR = '0') then
         s_Energy_Bin_227 <= s_Energy_Bin_227 +'1';
		 Energy_Bin_Rdy_227 <= '1';
		else
		 s_Energy_Bin_227 <= s_Energy_Bin_227;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_227 <= '0';
      end if;
    end if;
  end process  Energy_Bin_227;   
  
  Energy_Bin_228 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_228   <=  (others =>'0');
		Energy_Bin_Rdy_228 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E228_C1_L and PEAK_C1 <= s_E228_C1_H and Bin_OR = '0') then
         s_Energy_Bin_228 <= s_Energy_Bin_228 +'1';
		 Energy_Bin_Rdy_228 <= '1';
		else
		 s_Energy_Bin_228 <= s_Energy_Bin_228;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_228 <= '0';
      end if;
    end if;
  end process  Energy_Bin_228;   
  
  Energy_Bin_229 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_229   <=  (others =>'0');
		Energy_Bin_Rdy_229 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E229_C1_L and PEAK_C1 <= s_E229_C1_H and Bin_OR = '0') then
         s_Energy_Bin_229 <= s_Energy_Bin_229 +'1';
		 Energy_Bin_Rdy_229 <= '1';
		else
		 s_Energy_Bin_229 <= s_Energy_Bin_229;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_229 <= '0';
      end if;
    end if;
  end process  Energy_Bin_229;        
  
     Energy_Bin_230 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_230   <=  (others =>'0');
		Energy_Bin_Rdy_230 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E230_C1_L and PEAK_C1 <= s_E230_C1_H and Bin_OR = '0') then
         s_Energy_Bin_230 <= s_Energy_Bin_230 +'1';
		 Energy_Bin_Rdy_230 <= '1';
		else
		 s_Energy_Bin_230 <= s_Energy_Bin_230;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_230 <= '0';
      end if;
    end if;
  end process  Energy_Bin_230;    
  
  Energy_Bin_231 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_231   <=  (others =>'0');
		Energy_Bin_Rdy_231 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E231_C1_L and PEAK_C1 <= s_E231_C1_H and Bin_OR = '0') then
         s_Energy_Bin_231 <= s_Energy_Bin_231 +'1';
		 Energy_Bin_Rdy_231 <= '1';
		else
		 s_Energy_Bin_231 <= s_Energy_Bin_231;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_231 <= '0';
      end if;
    end if;
  end process  Energy_Bin_231;   
  
  Energy_Bin_232 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_232   <=  (others =>'0');
	    Energy_Bin_Rdy_232 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E232_C1_L and PEAK_C1 <= s_E232_C1_H and Bin_OR = '0') then
         s_Energy_Bin_232 <= s_Energy_Bin_232 +'1';
		 Energy_Bin_Rdy_232 <= '1';
		else
		 s_Energy_Bin_232 <= s_Energy_Bin_232;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_232 <= '0';
      end if;
    end if;
  end process  Energy_Bin_232;   
  
  Energy_Bin_233 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_233   <=  (others =>'0');
	    Energy_Bin_Rdy_233 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E233_C1_L and PEAK_C1 <= s_E233_C1_H and Bin_OR = '0') then
         s_Energy_Bin_233 <= s_Energy_Bin_233 +'1';
		 Energy_Bin_Rdy_233 <= '1';
		else
		 s_Energy_Bin_233 <= s_Energy_Bin_233;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_233 <= '0';
      end if;
    end if;
  end process  Energy_Bin_233;   
  
  Energy_Bin_234 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_234   <=  (others =>'0');
		Energy_Bin_Rdy_234 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E234_C1_L and PEAK_C1 <= s_E234_C1_H and Bin_OR = '0') then
         s_Energy_Bin_234 <= s_Energy_Bin_234 +'1';
		 Energy_Bin_Rdy_234 <= '1';
		else
		 s_Energy_Bin_234 <= s_Energy_Bin_234;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_234 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_234;   
 
 
  Energy_Bin_235 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_235   <=  (others =>'0');
		Energy_Bin_Rdy_235 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E235_C1_L and PEAK_C1 <= s_E235_C1_H and Bin_OR = '0') then
         s_Energy_Bin_235 <= s_Energy_Bin_235 +'1';
		 Energy_Bin_Rdy_235 <= '1';
		else
		 s_Energy_Bin_235 <= s_Energy_Bin_235;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_235 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_235;  
 
  
  Energy_Bin_236 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_236   <=  (others =>'0');
		Energy_Bin_Rdy_236 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E236_C1_L and PEAK_C1 <= s_E236_C1_H and Bin_OR = '0') then
         s_Energy_Bin_236 <= s_Energy_Bin_236 +'1';
		 Energy_Bin_Rdy_236 <= '1';
		else
		 s_Energy_Bin_236 <= s_Energy_Bin_236;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_236 <= '0';
      end if;
    end if;
  end process  Energy_Bin_236;   
  
 Energy_Bin_237 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_237   <=  (others =>'0');
		Energy_Bin_Rdy_237 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E237_C1_L and PEAK_C1 <= s_E237_C1_H and Bin_OR = '0') then
         s_Energy_Bin_237 <= s_Energy_Bin_237 +'1';
		 Energy_Bin_Rdy_237 <= '1';
		else
		 s_Energy_Bin_237 <= s_Energy_Bin_237;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_237 <= '0';
      end if;
    end if;
  end process  Energy_Bin_237;   
  
  Energy_Bin_238 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_238   <=  (others =>'0');
		Energy_Bin_Rdy_238 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E238_C1_L and PEAK_C1 <= s_E238_C1_H and Bin_OR = '0') then
         s_Energy_Bin_238 <= s_Energy_Bin_238 +'1';
		 Energy_Bin_Rdy_238 <= '1';
		else
		 s_Energy_Bin_238 <= s_Energy_Bin_238;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_238 <= '0';
      end if;
    end if;
  end process  Energy_Bin_238;   
  
  Energy_Bin_239 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_239   <=  (others =>'0');
		Energy_Bin_Rdy_239 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E239_C1_L and PEAK_C1 <= s_E239_C1_H and Bin_OR = '0') then
         s_Energy_Bin_239 <= s_Energy_Bin_239 +'1';
		 Energy_Bin_Rdy_239 <= '1';
		else
		 s_Energy_Bin_239 <= s_Energy_Bin_239;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_239 <= '0';
      end if;
    end if;
  end process  Energy_Bin_239;         
  
     Energy_Bin_240 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_240   <=  (others =>'0');
		Energy_Bin_Rdy_240 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E240_C1_L and PEAK_C1 <= s_E240_C1_H and Bin_OR = '0') then
         s_Energy_Bin_240 <= s_Energy_Bin_240 +'1';
		 Energy_Bin_Rdy_240 <= '1';
		else
		 s_Energy_Bin_240 <= s_Energy_Bin_240;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_240 <= '0';
      end if;
    end if;
  end process  Energy_Bin_240;    
  
  Energy_Bin_241 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_241   <=  (others =>'0');
		Energy_Bin_Rdy_241 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E241_C1_L and PEAK_C1 <= s_E241_C1_H and Bin_OR = '0') then
         s_Energy_Bin_241 <= s_Energy_Bin_241 +'1';
		 Energy_Bin_Rdy_241 <= '1';
		else
		 s_Energy_Bin_241 <= s_Energy_Bin_241;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_241 <= '0';
      end if;
    end if;
  end process  Energy_Bin_241;   
  
  Energy_Bin_242 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_242   <=  (others =>'0');
	    Energy_Bin_Rdy_242 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E242_C1_L and PEAK_C1 <= s_E242_C1_H and Bin_OR = '0') then
         s_Energy_Bin_242 <= s_Energy_Bin_242 +'1';
		 Energy_Bin_Rdy_242 <= '1';
		else
		 s_Energy_Bin_242 <= s_Energy_Bin_242;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_242 <= '0';
      end if;
    end if;
  end process  Energy_Bin_242;   
  
  Energy_Bin_243 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_243   <=  (others =>'0');
	    Energy_Bin_Rdy_243 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E243_C1_L and PEAK_C1 <= s_E243_C1_H and Bin_OR = '0') then
         s_Energy_Bin_243 <= s_Energy_Bin_243 +'1';
		 Energy_Bin_Rdy_243 <= '1';
		else
		 s_Energy_Bin_243 <= s_Energy_Bin_243;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_243 <= '0';
      end if;
    end if;
  end process  Energy_Bin_243;   
  
  Energy_Bin_244 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_244   <=  (others =>'0');
		Energy_Bin_Rdy_244 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E244_C1_L and PEAK_C1 <= s_E244_C1_H and Bin_OR = '0') then
         s_Energy_Bin_244 <= s_Energy_Bin_244 +'1';
		 Energy_Bin_Rdy_244 <= '1';
		else
		 s_Energy_Bin_244 <= s_Energy_Bin_244;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_244 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_244;   
 
 
  Energy_Bin_245 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_245   <=  (others =>'0');
		Energy_Bin_Rdy_245 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E245_C1_L and PEAK_C1 <= s_E245_C1_H and Bin_OR = '0') then
         s_Energy_Bin_245 <= s_Energy_Bin_245 +'1';
		 Energy_Bin_Rdy_245 <= '1';
		else
		 s_Energy_Bin_245 <= s_Energy_Bin_245;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_245 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_245;  
 
  
  Energy_Bin_246 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_246   <=  (others =>'0');
		Energy_Bin_Rdy_246 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E246_C1_L and PEAK_C1 <= s_E246_C1_H and Bin_OR = '0') then
         s_Energy_Bin_246 <= s_Energy_Bin_246 +'1';
		 Energy_Bin_Rdy_246 <= '1';
		else
		 s_Energy_Bin_246 <= s_Energy_Bin_246;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_246 <= '0';
      end if;
    end if;
  end process  Energy_Bin_246;   
  
 Energy_Bin_247 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_247   <=  (others =>'0');
		Energy_Bin_Rdy_247 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E247_C1_L and PEAK_C1 <= s_E247_C1_H and Bin_OR = '0') then
         s_Energy_Bin_247 <= s_Energy_Bin_247 +'1';
		 Energy_Bin_Rdy_247 <= '1';
		else
		 s_Energy_Bin_247 <= s_Energy_Bin_247;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_247 <= '0';
      end if;
    end if;
  end process  Energy_Bin_247;   
  
  Energy_Bin_248 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_248   <=  (others =>'0');
		Energy_Bin_Rdy_248 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E248_C1_L and PEAK_C1 <= s_E248_C1_H and Bin_OR = '0') then
         s_Energy_Bin_248 <= s_Energy_Bin_248 +'1';
		 Energy_Bin_Rdy_248 <= '1';
		else
		 s_Energy_Bin_248 <= s_Energy_Bin_248;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_248 <= '0';
      end if;
    end if;
  end process  Energy_Bin_248;   
  
  Energy_Bin_249 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_249   <=  (others =>'0');
		Energy_Bin_Rdy_249 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E249_C1_L and PEAK_C1 <= s_E249_C1_H and Bin_OR = '0') then
         s_Energy_Bin_249 <= s_Energy_Bin_249 +'1';
		 Energy_Bin_Rdy_249 <= '1';
		else
		 s_Energy_Bin_249 <= s_Energy_Bin_249;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_249 <= '0';
      end if;
    end if;
  end process  Energy_Bin_249;          
  
  
     Energy_Bin_250 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_250   <=  (others =>'0');
		Energy_Bin_Rdy_250 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E250_C1_L and PEAK_C1 <= s_E250_C1_H and Bin_OR = '0') then
         s_Energy_Bin_250 <= s_Energy_Bin_250 +'1';
		 Energy_Bin_Rdy_250 <= '1';
		else
		 s_Energy_Bin_250 <= s_Energy_Bin_250;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_250 <= '0';
      end if;
    end if;
  end process  Energy_Bin_250;    
  
  Energy_Bin_251 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_251   <=  (others =>'0');
		Energy_Bin_Rdy_251 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E251_C1_L and PEAK_C1 <= s_E251_C1_H and Bin_OR = '0') then
         s_Energy_Bin_251 <= s_Energy_Bin_251 +'1';
		 Energy_Bin_Rdy_251 <= '1';
		else
		 s_Energy_Bin_251 <= s_Energy_Bin_251;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_251 <= '0';
      end if;
    end if;
  end process  Energy_Bin_251;   
  
  Energy_Bin_252 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_252   <=  (others =>'0');
	    Energy_Bin_Rdy_252 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E252_C1_L and PEAK_C1 <= s_E252_C1_H and Bin_OR = '0') then
         s_Energy_Bin_252 <= s_Energy_Bin_252 +'1';
		 Energy_Bin_Rdy_252 <= '1';
		else
		 s_Energy_Bin_252 <= s_Energy_Bin_252;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_252 <= '0';
      end if;
    end if;
  end process  Energy_Bin_252;   
  
  Energy_Bin_253 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_253   <=  (others =>'0');
	    Energy_Bin_Rdy_253 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E253_C1_L and PEAK_C1 <= s_E253_C1_H and Bin_OR = '0') then
         s_Energy_Bin_253 <= s_Energy_Bin_253 +'1';
		 Energy_Bin_Rdy_253 <= '1';
		else
		 s_Energy_Bin_253 <= s_Energy_Bin_253;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_253 <= '0';
      end if;
    end if;
  end process  Energy_Bin_253;   
  
  Energy_Bin_254 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_254   <=  (others =>'0');
		Energy_Bin_Rdy_254 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E254_C1_L and PEAK_C1 <= s_E254_C1_H and Bin_OR = '0') then
         s_Energy_Bin_254 <= s_Energy_Bin_254 +'1';
		 Energy_Bin_Rdy_254 <= '1';
		else
		 s_Energy_Bin_254 <= s_Energy_Bin_254;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_254 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_254;   
 
 
  Energy_Bin_255 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_255   <=  (others =>'0');
		Energy_Bin_Rdy_255 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E255_C1_L and PEAK_C1 <= s_E255_C1_H and Bin_OR = '0') then
         s_Energy_Bin_255 <= s_Energy_Bin_255 +'1';
		 Energy_Bin_Rdy_255 <= '1';
		else
		 s_Energy_Bin_255 <= s_Energy_Bin_255;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_255 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_255;  
 
  
  Energy_Bin_256 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_256   <=  (others =>'0');
		Energy_Bin_Rdy_256 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E256_C1_L and PEAK_C1 <= s_E256_C1_H and Bin_OR = '0') then
         s_Energy_Bin_256 <= s_Energy_Bin_256 +'1';
		 Energy_Bin_Rdy_256 <= '1';
		else
		 s_Energy_Bin_256 <= s_Energy_Bin_256;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_256 <= '0';
      end if;
    end if;
  end process  Energy_Bin_256;   
  
 Energy_Bin_257 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_257   <=  (others =>'0');
		Energy_Bin_Rdy_257 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E257_C1_L and PEAK_C1 <= s_E257_C1_H and Bin_OR = '0') then
         s_Energy_Bin_257 <= s_Energy_Bin_257 +'1';
		 Energy_Bin_Rdy_257 <= '1';
		else
		 s_Energy_Bin_257 <= s_Energy_Bin_257;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_257 <= '0';
      end if;
    end if;
  end process  Energy_Bin_257;   
  
  Energy_Bin_258 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_258   <=  (others =>'0');
		Energy_Bin_Rdy_258 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E258_C1_L and PEAK_C1 <= s_E258_C1_H and Bin_OR = '0') then
         s_Energy_Bin_258 <= s_Energy_Bin_258 +'1';
		 Energy_Bin_Rdy_258 <= '1';
		else
		 s_Energy_Bin_258 <= s_Energy_Bin_258;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_258 <= '0';
      end if;
    end if;
  end process  Energy_Bin_258;   
  
  Energy_Bin_259 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_259   <=  (others =>'0');
		Energy_Bin_Rdy_259 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E259_C1_L and PEAK_C1 <= s_E259_C1_H and Bin_OR = '0') then
         s_Energy_Bin_259 <= s_Energy_Bin_259 +'1';
		 Energy_Bin_Rdy_259 <= '1';
		else
		 s_Energy_Bin_259 <= s_Energy_Bin_259;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_259 <= '0';
      end if;
    end if;
  end process  Energy_Bin_259;           
  
     Energy_Bin_260 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_260   <=  (others =>'0');
		Energy_Bin_Rdy_260 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E260_C1_L and PEAK_C1 <= s_E260_C1_H and Bin_OR = '0') then
         s_Energy_Bin_260 <= s_Energy_Bin_260 +'1';
		 Energy_Bin_Rdy_260 <= '1';
		else
		 s_Energy_Bin_260 <= s_Energy_Bin_260;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_260 <= '0';
      end if;
    end if;
  end process  Energy_Bin_260;    
  
  Energy_Bin_261 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_261   <=  (others =>'0');
		Energy_Bin_Rdy_261 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E261_C1_L and PEAK_C1 <= s_E261_C1_H and Bin_OR = '0') then
         s_Energy_Bin_261 <= s_Energy_Bin_261 +'1';
		 Energy_Bin_Rdy_261 <= '1';
		else
		 s_Energy_Bin_261 <= s_Energy_Bin_261;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_261 <= '0';
      end if;
    end if;
  end process  Energy_Bin_261;   
  
  Energy_Bin_262 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_262   <=  (others =>'0');
	    Energy_Bin_Rdy_262 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E262_C1_L and PEAK_C1 <= s_E262_C1_H and Bin_OR = '0') then
         s_Energy_Bin_262 <= s_Energy_Bin_262 +'1';
		 Energy_Bin_Rdy_262 <= '1';
		else
		 s_Energy_Bin_262 <= s_Energy_Bin_262;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_262 <= '0';
      end if;
    end if;
  end process  Energy_Bin_262;   
  
  Energy_Bin_263 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_263   <=  (others =>'0');
	    Energy_Bin_Rdy_263 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E263_C1_L and PEAK_C1 <= s_E263_C1_H and Bin_OR = '0') then
         s_Energy_Bin_263 <= s_Energy_Bin_263 +'1';
		 Energy_Bin_Rdy_263 <= '1';
		else
		 s_Energy_Bin_263 <= s_Energy_Bin_263;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_263 <= '0';
      end if;
    end if;
  end process  Energy_Bin_263;   
  
  Energy_Bin_264 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_264   <=  (others =>'0');
		Energy_Bin_Rdy_264 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E264_C1_L and PEAK_C1 <= s_E264_C1_H and Bin_OR = '0') then
         s_Energy_Bin_264 <= s_Energy_Bin_264 +'1';
		 Energy_Bin_Rdy_264 <= '1';
		else
		 s_Energy_Bin_264 <= s_Energy_Bin_264;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_264 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_264;   
 
 
  Energy_Bin_265 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_265   <=  (others =>'0');
		Energy_Bin_Rdy_265 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E265_C1_L and PEAK_C1 <= s_E265_C1_H and Bin_OR = '0') then
         s_Energy_Bin_265 <= s_Energy_Bin_265 +'1';
		 Energy_Bin_Rdy_265 <= '1';
		else
		 s_Energy_Bin_265 <= s_Energy_Bin_265;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_265 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_265;  
 
  
  Energy_Bin_266 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_266   <=  (others =>'0');
		Energy_Bin_Rdy_266 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E266_C1_L and PEAK_C1 <= s_E266_C1_H and Bin_OR = '0') then
         s_Energy_Bin_266 <= s_Energy_Bin_266 +'1';
		 Energy_Bin_Rdy_266 <= '1';
		else
		 s_Energy_Bin_266 <= s_Energy_Bin_266;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_266 <= '0';
      end if;
    end if;
  end process  Energy_Bin_266;   
  
 Energy_Bin_267 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_267   <=  (others =>'0');
		Energy_Bin_Rdy_267 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E267_C1_L and PEAK_C1 <= s_E267_C1_H and Bin_OR = '0') then
         s_Energy_Bin_267 <= s_Energy_Bin_267 +'1';
		 Energy_Bin_Rdy_267 <= '1';
		else
		 s_Energy_Bin_267 <= s_Energy_Bin_267;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_267 <= '0';
      end if;
    end if;
  end process  Energy_Bin_267;   
  
  Energy_Bin_268 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_268   <=  (others =>'0');
		Energy_Bin_Rdy_268 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E268_C1_L and PEAK_C1 <= s_E268_C1_H and Bin_OR = '0') then
         s_Energy_Bin_268 <= s_Energy_Bin_268 +'1';
		 Energy_Bin_Rdy_268 <= '1';
		else
		 s_Energy_Bin_268 <= s_Energy_Bin_268;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_268 <= '0';
      end if;
    end if;
  end process  Energy_Bin_268;   
  
  Energy_Bin_269 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_269   <=  (others =>'0');
		Energy_Bin_Rdy_269 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E269_C1_L and PEAK_C1 <= s_E269_C1_H and Bin_OR = '0') then
         s_Energy_Bin_269 <= s_Energy_Bin_269 +'1';
		 Energy_Bin_Rdy_269 <= '1';
		else
		 s_Energy_Bin_269 <= s_Energy_Bin_269;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_269 <= '0';
      end if;
    end if;
  end process  Energy_Bin_269;         
  
     Energy_Bin_270 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_270   <=  (others =>'0');
		Energy_Bin_Rdy_270 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E270_C1_L and PEAK_C1 <= s_E270_C1_H and Bin_OR = '0') then
         s_Energy_Bin_270 <= s_Energy_Bin_270 +'1';
		 Energy_Bin_Rdy_270 <= '1';
		else
		 s_Energy_Bin_270 <= s_Energy_Bin_270;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_270 <= '0';
      end if;
    end if;
  end process  Energy_Bin_270;    
  
  Energy_Bin_271 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_271   <=  (others =>'0');
		Energy_Bin_Rdy_271 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E271_C1_L and PEAK_C1 <= s_E271_C1_H and Bin_OR = '0') then
         s_Energy_Bin_271 <= s_Energy_Bin_271 +'1';
		 Energy_Bin_Rdy_271 <= '1';
		else
		 s_Energy_Bin_271 <= s_Energy_Bin_271;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_271 <= '0';
      end if;
    end if;
  end process  Energy_Bin_271;   
  
  Energy_Bin_272 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_272   <=  (others =>'0');
	    Energy_Bin_Rdy_272 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E272_C1_L and PEAK_C1 <= s_E272_C1_H and Bin_OR = '0') then
         s_Energy_Bin_272 <= s_Energy_Bin_272 +'1';
		 Energy_Bin_Rdy_272 <= '1';
		else
		 s_Energy_Bin_272 <= s_Energy_Bin_272;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_272 <= '0';
      end if;
    end if;
  end process  Energy_Bin_272;   
  
  Energy_Bin_273 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_273   <=  (others =>'0');
	    Energy_Bin_Rdy_273 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E273_C1_L and PEAK_C1 <= s_E273_C1_H and Bin_OR = '0') then
         s_Energy_Bin_273 <= s_Energy_Bin_273 +'1';
		 Energy_Bin_Rdy_273 <= '1';
		else
		 s_Energy_Bin_273 <= s_Energy_Bin_273;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_273 <= '0';
      end if;
    end if;
  end process  Energy_Bin_273;   
  
  Energy_Bin_274 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_274   <=  (others =>'0');
		Energy_Bin_Rdy_274 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E274_C1_L and PEAK_C1 <= s_E274_C1_H and Bin_OR = '0') then
         s_Energy_Bin_274 <= s_Energy_Bin_274 +'1';
		 Energy_Bin_Rdy_274 <= '1';
		else
		 s_Energy_Bin_274 <= s_Energy_Bin_274;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_274 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_274;   
 
 
  Energy_Bin_275 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_275   <=  (others =>'0');
		Energy_Bin_Rdy_275 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E275_C1_L and PEAK_C1 <= s_E275_C1_H and Bin_OR = '0') then
         s_Energy_Bin_275 <= s_Energy_Bin_275 +'1';
		 Energy_Bin_Rdy_275 <= '1';
		else
		 s_Energy_Bin_275 <= s_Energy_Bin_275;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_275 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_275;  
 
  
  Energy_Bin_276 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_276   <=  (others =>'0');
		Energy_Bin_Rdy_276 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E276_C1_L and PEAK_C1 <= s_E276_C1_H and Bin_OR = '0') then
         s_Energy_Bin_276 <= s_Energy_Bin_276 +'1';
		 Energy_Bin_Rdy_276 <= '1';
		else
		 s_Energy_Bin_276 <= s_Energy_Bin_276;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_276 <= '0';
      end if;
    end if;
  end process  Energy_Bin_276;   
  
 Energy_Bin_277 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_277   <=  (others =>'0');
		Energy_Bin_Rdy_277 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E277_C1_L and PEAK_C1 <= s_E277_C1_H and Bin_OR = '0') then
         s_Energy_Bin_277 <= s_Energy_Bin_277 +'1';
		 Energy_Bin_Rdy_277 <= '1';
		else
		 s_Energy_Bin_277 <= s_Energy_Bin_277;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_277 <= '0';
      end if;
    end if;
  end process  Energy_Bin_277;   
  
  Energy_Bin_278 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_278   <=  (others =>'0');
		Energy_Bin_Rdy_278 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E278_C1_L and PEAK_C1 <= s_E278_C1_H and Bin_OR = '0') then
         s_Energy_Bin_278 <= s_Energy_Bin_278 +'1';
		 Energy_Bin_Rdy_278 <= '1';
		else
		 s_Energy_Bin_278 <= s_Energy_Bin_278;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_278 <= '0';
      end if;
    end if;
  end process  Energy_Bin_278;   
  
  Energy_Bin_279 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_279   <=  (others =>'0');
		Energy_Bin_Rdy_279 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E279_C1_L and PEAK_C1 <= s_E279_C1_H and Bin_OR = '0') then
         s_Energy_Bin_279 <= s_Energy_Bin_279 +'1';
		 Energy_Bin_Rdy_279 <= '1';
		else
		 s_Energy_Bin_279 <= s_Energy_Bin_279;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_279 <= '0';
      end if;
    end if;
  end process  Energy_Bin_279;       
  
     Energy_Bin_280 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_280   <=  (others =>'0');
		Energy_Bin_Rdy_280 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E280_C1_L and PEAK_C1 <= s_E280_C1_H and Bin_OR = '0') then
         s_Energy_Bin_280 <= s_Energy_Bin_280 +'1';
		 Energy_Bin_Rdy_280 <= '1';
		else
		 s_Energy_Bin_280 <= s_Energy_Bin_280;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_280 <= '0';
      end if;
    end if;
  end process  Energy_Bin_280;    
  
  Energy_Bin_281 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_281   <=  (others =>'0');
		Energy_Bin_Rdy_281 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E281_C1_L and PEAK_C1 <= s_E281_C1_H and Bin_OR = '0') then
         s_Energy_Bin_281 <= s_Energy_Bin_281 +'1';
		 Energy_Bin_Rdy_281 <= '1';
		else
		 s_Energy_Bin_281 <= s_Energy_Bin_281;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_281 <= '0';
      end if;
    end if;
  end process  Energy_Bin_281;   
  
  Energy_Bin_282 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_282   <=  (others =>'0');
	    Energy_Bin_Rdy_282 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E282_C1_L and PEAK_C1 <= s_E282_C1_H and Bin_OR = '0') then
         s_Energy_Bin_282 <= s_Energy_Bin_282 +'1';
		 Energy_Bin_Rdy_282 <= '1';
		else
		 s_Energy_Bin_282 <= s_Energy_Bin_282;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_282 <= '0';
      end if;
    end if;
  end process  Energy_Bin_282;   
  
  Energy_Bin_283 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_283   <=  (others =>'0');
	    Energy_Bin_Rdy_283 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E283_C1_L and PEAK_C1 <= s_E283_C1_H and Bin_OR = '0') then
         s_Energy_Bin_283 <= s_Energy_Bin_283 +'1';
		 Energy_Bin_Rdy_283 <= '1';
		else
		 s_Energy_Bin_283 <= s_Energy_Bin_283;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_283 <= '0';
      end if;
    end if;
  end process  Energy_Bin_283;   
  
  Energy_Bin_284 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_284   <=  (others =>'0');
		Energy_Bin_Rdy_284 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E284_C1_L and PEAK_C1 <= s_E284_C1_H and Bin_OR = '0') then
         s_Energy_Bin_284 <= s_Energy_Bin_284 +'1';
		 Energy_Bin_Rdy_284 <= '1';
		else
		 s_Energy_Bin_284 <= s_Energy_Bin_284;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_284 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_284;   
 
 
  Energy_Bin_285 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_285   <=  (others =>'0');
		Energy_Bin_Rdy_285 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E285_C1_L and PEAK_C1 <= s_E285_C1_H and Bin_OR = '0') then
         s_Energy_Bin_285 <= s_Energy_Bin_285 +'1';
		 Energy_Bin_Rdy_285 <= '1';
		else
		 s_Energy_Bin_285 <= s_Energy_Bin_285;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_285 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_285;  
 
  
  Energy_Bin_286 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_286   <=  (others =>'0');
		Energy_Bin_Rdy_286 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E286_C1_L and PEAK_C1 <= s_E286_C1_H and Bin_OR = '0') then
         s_Energy_Bin_286 <= s_Energy_Bin_286 +'1';
		 Energy_Bin_Rdy_286 <= '1';
		else
		 s_Energy_Bin_286 <= s_Energy_Bin_286;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_286 <= '0';
      end if;
    end if;
  end process  Energy_Bin_286;   
  
 Energy_Bin_287 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_287   <=  (others =>'0');
		Energy_Bin_Rdy_287 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E287_C1_L and PEAK_C1 <= s_E287_C1_H and Bin_OR = '0') then
         s_Energy_Bin_287 <= s_Energy_Bin_287 +'1';
		 Energy_Bin_Rdy_287 <= '1';
		else
		 s_Energy_Bin_287 <= s_Energy_Bin_287;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_287 <= '0';
      end if;
    end if;
  end process  Energy_Bin_287;   
  
  Energy_Bin_288 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_288   <=  (others =>'0');
		Energy_Bin_Rdy_288 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E288_C1_L and PEAK_C1 <= s_E288_C1_H and Bin_OR = '0') then
         s_Energy_Bin_288 <= s_Energy_Bin_288 +'1';
		 Energy_Bin_Rdy_288 <= '1';
		else
		 s_Energy_Bin_288 <= s_Energy_Bin_288;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_288 <= '0';
      end if;
    end if;
  end process  Energy_Bin_288;   
  
  Energy_Bin_289 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_289   <=  (others =>'0');
		Energy_Bin_Rdy_289 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E289_C1_L and PEAK_C1 <= s_E289_C1_H and Bin_OR = '0') then
         s_Energy_Bin_289 <= s_Energy_Bin_289 +'1';
		 Energy_Bin_Rdy_289 <= '1';
		else
		 s_Energy_Bin_289 <= s_Energy_Bin_289;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_289 <= '0';
      end if;
    end if;
  end process  Energy_Bin_289;      
  
     Energy_Bin_290 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_290   <=  (others =>'0');
		Energy_Bin_Rdy_290 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E290_C1_L and PEAK_C1 <= s_E290_C1_H and Bin_OR = '0') then
         s_Energy_Bin_290 <= s_Energy_Bin_290 +'1';
		 Energy_Bin_Rdy_290 <= '1';
		else
		 s_Energy_Bin_290 <= s_Energy_Bin_290;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_290 <= '0';
      end if;
    end if;
  end process  Energy_Bin_290;    
  
  Energy_Bin_291 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_291   <=  (others =>'0');
		Energy_Bin_Rdy_291 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E291_C1_L and PEAK_C1 <= s_E291_C1_H and Bin_OR = '0') then
         s_Energy_Bin_291 <= s_Energy_Bin_291 +'1';
		 Energy_Bin_Rdy_291 <= '1';
		else
		 s_Energy_Bin_291 <= s_Energy_Bin_291;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_291 <= '0';
      end if;
    end if;
  end process  Energy_Bin_291;   
  
  Energy_Bin_292 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_292   <=  (others =>'0');
	    Energy_Bin_Rdy_292 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E292_C1_L and PEAK_C1 <= s_E292_C1_H and Bin_OR = '0') then
         s_Energy_Bin_292 <= s_Energy_Bin_292 +'1';
		 Energy_Bin_Rdy_292 <= '1';
		else
		 s_Energy_Bin_292 <= s_Energy_Bin_292;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_292 <= '0';
      end if;
    end if;
  end process  Energy_Bin_292;   
  
  Energy_Bin_293 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_293   <=  (others =>'0');
	    Energy_Bin_Rdy_293 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E293_C1_L and PEAK_C1 <= s_E293_C1_H and Bin_OR = '0') then
         s_Energy_Bin_293 <= s_Energy_Bin_293 +'1';
		 Energy_Bin_Rdy_293 <= '1';
		else
		 s_Energy_Bin_293 <= s_Energy_Bin_293;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_293 <= '0';
      end if;
    end if;
  end process  Energy_Bin_293;   
  
  Energy_Bin_294 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_294   <=  (others =>'0');
		Energy_Bin_Rdy_294 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E294_C1_L and PEAK_C1 <= s_E294_C1_H and Bin_OR = '0') then
         s_Energy_Bin_294 <= s_Energy_Bin_294 +'1';
		 Energy_Bin_Rdy_294 <= '1';
		else
		 s_Energy_Bin_294 <= s_Energy_Bin_294;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_294 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_294;   
 
 
  Energy_Bin_295 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_295   <=  (others =>'0');
		Energy_Bin_Rdy_295 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E295_C1_L and PEAK_C1 <= s_E295_C1_H and Bin_OR = '0') then
         s_Energy_Bin_295 <= s_Energy_Bin_295 +'1';
		 Energy_Bin_Rdy_295 <= '1';
		else
		 s_Energy_Bin_295 <= s_Energy_Bin_295;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_295 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_295;  
 
  
  Energy_Bin_296 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_296   <=  (others =>'0');
		Energy_Bin_Rdy_296 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E296_C1_L and PEAK_C1 <= s_E296_C1_H and Bin_OR = '0') then
         s_Energy_Bin_296 <= s_Energy_Bin_296 +'1';
		 Energy_Bin_Rdy_296 <= '1';
		else
		 s_Energy_Bin_296 <= s_Energy_Bin_296;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_296 <= '0';
      end if;
    end if;
  end process  Energy_Bin_296;   
  
 Energy_Bin_297 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_297   <=  (others =>'0');
		Energy_Bin_Rdy_297 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E297_C1_L and PEAK_C1 <= s_E297_C1_H and Bin_OR = '0') then
         s_Energy_Bin_297 <= s_Energy_Bin_297 +'1';
		 Energy_Bin_Rdy_297 <= '1';
		else
		 s_Energy_Bin_297 <= s_Energy_Bin_297;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_297 <= '0';
      end if;
    end if;
  end process  Energy_Bin_297;   
  
  Energy_Bin_298 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_298   <=  (others =>'0');
		Energy_Bin_Rdy_298 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E298_C1_L and PEAK_C1 <= s_E298_C1_H and Bin_OR = '0') then
         s_Energy_Bin_298 <= s_Energy_Bin_298 +'1';
		 Energy_Bin_Rdy_298 <= '1';
		else
		 s_Energy_Bin_298 <= s_Energy_Bin_298;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_298 <= '0';
      end if;
    end if;
  end process  Energy_Bin_298;   
  
  Energy_Bin_299 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_299   <=  (others =>'0');
		Energy_Bin_Rdy_299 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E299_C1_L and PEAK_C1 <= s_E299_C1_H and Bin_OR = '0') then
         s_Energy_Bin_299 <= s_Energy_Bin_299 +'1';
		 Energy_Bin_Rdy_299 <= '1';
		else
		 s_Energy_Bin_299 <= s_Energy_Bin_299;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_299 <= '0';
      end if;
    end if;
  end process  Energy_Bin_299;      

     Energy_Bin_300 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_300   <=  (others =>'0');
		Energy_Bin_Rdy_300 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E300_C1_L and PEAK_C1 <= s_E300_C1_H and Bin_OR = '0') then
         s_Energy_Bin_300 <= s_Energy_Bin_300 +'1';
		 Energy_Bin_Rdy_300 <= '1';
		else
		 s_Energy_Bin_300 <= s_Energy_Bin_300;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_300 <= '0';
      end if;
    end if;
  end process  Energy_Bin_300;    
  
  Energy_Bin_301 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_301   <=  (others =>'0');
		Energy_Bin_Rdy_301 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E301_C1_L and PEAK_C1 <= s_E301_C1_H and Bin_OR = '0') then
         s_Energy_Bin_301 <= s_Energy_Bin_301 +'1';
		 Energy_Bin_Rdy_301 <= '1';
		else
		 s_Energy_Bin_301 <= s_Energy_Bin_301;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_301 <= '0';
      end if;
    end if;
  end process  Energy_Bin_301;   
  
  Energy_Bin_302 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_302   <=  (others =>'0');
	    Energy_Bin_Rdy_302 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E302_C1_L and PEAK_C1 <= s_E302_C1_H and Bin_OR = '0') then
         s_Energy_Bin_302 <= s_Energy_Bin_302 +'1';
		 Energy_Bin_Rdy_302 <= '1';
		else
		 s_Energy_Bin_302 <= s_Energy_Bin_302;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_302 <= '0';
      end if;
    end if;
  end process  Energy_Bin_302;   
  
  Energy_Bin_303 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_303   <=  (others =>'0');
	    Energy_Bin_Rdy_303 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E303_C1_L and PEAK_C1 <= s_E303_C1_H and Bin_OR = '0') then
         s_Energy_Bin_303 <= s_Energy_Bin_303 +'1';
		 Energy_Bin_Rdy_303 <= '1';
		else
		 s_Energy_Bin_303 <= s_Energy_Bin_303;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_303 <= '0';
      end if;
    end if;
  end process  Energy_Bin_303;   
  
  Energy_Bin_304 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_304   <=  (others =>'0');
		Energy_Bin_Rdy_304 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E304_C1_L and PEAK_C1 <= s_E304_C1_H and Bin_OR = '0') then
         s_Energy_Bin_304 <= s_Energy_Bin_304 +'1';
		 Energy_Bin_Rdy_304 <= '1';
		else
		 s_Energy_Bin_304 <= s_Energy_Bin_304;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_304 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_304;   
 
 
  Energy_Bin_305 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_305   <=  (others =>'0');
		Energy_Bin_Rdy_305 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E305_C1_L and PEAK_C1 <= s_E305_C1_H and Bin_OR = '0') then
         s_Energy_Bin_305 <= s_Energy_Bin_305 +'1';
		 Energy_Bin_Rdy_305 <= '1';
		else
		 s_Energy_Bin_305 <= s_Energy_Bin_305;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_305 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_305;  
 
  
  Energy_Bin_306 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_306   <=  (others =>'0');
		Energy_Bin_Rdy_306 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E306_C1_L and PEAK_C1 <= s_E306_C1_H and Bin_OR = '0') then
         s_Energy_Bin_306 <= s_Energy_Bin_306 +'1';
		 Energy_Bin_Rdy_306 <= '1';
		else
		 s_Energy_Bin_306 <= s_Energy_Bin_306;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_306 <= '0';
      end if;
    end if;
  end process  Energy_Bin_306;   
  
 Energy_Bin_307 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_307   <=  (others =>'0');
		Energy_Bin_Rdy_307 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E307_C1_L and PEAK_C1 <= s_E307_C1_H and Bin_OR = '0') then
         s_Energy_Bin_307 <= s_Energy_Bin_307 +'1';
		 Energy_Bin_Rdy_307 <= '1';
		else
		 s_Energy_Bin_307 <= s_Energy_Bin_307;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_307 <= '0';
      end if;
    end if;
  end process  Energy_Bin_307;   
  
  Energy_Bin_308 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_308   <=  (others =>'0');
		Energy_Bin_Rdy_308 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E308_C1_L and PEAK_C1 <= s_E308_C1_H and Bin_OR = '0') then
         s_Energy_Bin_308 <= s_Energy_Bin_308 +'1';
		 Energy_Bin_Rdy_308 <= '1';
		else
		 s_Energy_Bin_308 <= s_Energy_Bin_308;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_308 <= '0';
      end if;
    end if;
  end process  Energy_Bin_308;   
  
  Energy_Bin_309 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_309   <=  (others =>'0');
		Energy_Bin_Rdy_309 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E309_C1_L and PEAK_C1 <= s_E309_C1_H and Bin_OR = '0') then
         s_Energy_Bin_309 <= s_Energy_Bin_309 +'1';
		 Energy_Bin_Rdy_309 <= '1';
		else
		 s_Energy_Bin_309 <= s_Energy_Bin_309;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_309 <= '0';
      end if;
    end if;
  end process  Energy_Bin_309;      
  
     Energy_Bin_310 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_310   <=  (others =>'0');
		Energy_Bin_Rdy_310 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E310_C1_L and PEAK_C1 <= s_E310_C1_H and Bin_OR = '0') then
         s_Energy_Bin_310 <= s_Energy_Bin_310 +'1';
		 Energy_Bin_Rdy_310 <= '1';
		else
		 s_Energy_Bin_310 <= s_Energy_Bin_310;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_310 <= '0';
      end if;
    end if;
  end process  Energy_Bin_310;    
  
  Energy_Bin_311 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_311   <=  (others =>'0');
		Energy_Bin_Rdy_311 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E311_C1_L and PEAK_C1 <= s_E311_C1_H and Bin_OR = '0') then
         s_Energy_Bin_311 <= s_Energy_Bin_311 +'1';
		 Energy_Bin_Rdy_311 <= '1';
		else
		 s_Energy_Bin_311 <= s_Energy_Bin_311;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_311 <= '0';
      end if;
    end if;
  end process  Energy_Bin_311;   
  
  Energy_Bin_312 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_312   <=  (others =>'0');
	    Energy_Bin_Rdy_312 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E312_C1_L and PEAK_C1 <= s_E312_C1_H and Bin_OR = '0') then
         s_Energy_Bin_312 <= s_Energy_Bin_312 +'1';
		 Energy_Bin_Rdy_312 <= '1';
		else
		 s_Energy_Bin_312 <= s_Energy_Bin_312;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_312 <= '0';
      end if;
    end if;
  end process  Energy_Bin_312;   
  
  Energy_Bin_313 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_313   <=  (others =>'0');
	    Energy_Bin_Rdy_313 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E313_C1_L and PEAK_C1 <= s_E313_C1_H and Bin_OR = '0') then
         s_Energy_Bin_313 <= s_Energy_Bin_313 +'1';
		 Energy_Bin_Rdy_313 <= '1';
		else
		 s_Energy_Bin_313 <= s_Energy_Bin_313;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_313 <= '0';
      end if;
    end if;
  end process  Energy_Bin_313;   
  
  Energy_Bin_314 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_314   <=  (others =>'0');
		Energy_Bin_Rdy_314 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E314_C1_L and PEAK_C1 <= s_E314_C1_H and Bin_OR = '0') then
         s_Energy_Bin_314 <= s_Energy_Bin_314 +'1';
		 Energy_Bin_Rdy_314 <= '1';
		else
		 s_Energy_Bin_314 <= s_Energy_Bin_314;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_314 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_314;   
 
 
  Energy_Bin_315 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_315   <=  (others =>'0');
		Energy_Bin_Rdy_315 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E315_C1_L and PEAK_C1 <= s_E315_C1_H and Bin_OR = '0') then
         s_Energy_Bin_315 <= s_Energy_Bin_315 +'1';
		 Energy_Bin_Rdy_315 <= '1';
		else
		 s_Energy_Bin_315 <= s_Energy_Bin_315;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_315 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_315;  
 
  
  Energy_Bin_316 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_316   <=  (others =>'0');
		Energy_Bin_Rdy_316 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E316_C1_L and PEAK_C1 <= s_E316_C1_H and Bin_OR = '0') then
         s_Energy_Bin_316 <= s_Energy_Bin_316 +'1';
		 Energy_Bin_Rdy_316 <= '1';
		else
		 s_Energy_Bin_316 <= s_Energy_Bin_316;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_316 <= '0';
      end if;
    end if;
  end process  Energy_Bin_316;   
  
 Energy_Bin_317 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_317   <=  (others =>'0');
		Energy_Bin_Rdy_317 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E317_C1_L and PEAK_C1 <= s_E317_C1_H and Bin_OR = '0') then
         s_Energy_Bin_317 <= s_Energy_Bin_317 +'1';
		 Energy_Bin_Rdy_317 <= '1';
		else
		 s_Energy_Bin_317 <= s_Energy_Bin_317;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_317 <= '0';
      end if;
    end if;
  end process  Energy_Bin_317;   
  
  Energy_Bin_318 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_318   <=  (others =>'0');
		Energy_Bin_Rdy_318 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E318_C1_L and PEAK_C1 <= s_E318_C1_H and Bin_OR = '0') then
         s_Energy_Bin_318 <= s_Energy_Bin_318 +'1';
		 Energy_Bin_Rdy_318 <= '1';
		else
		 s_Energy_Bin_318 <= s_Energy_Bin_318;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_318 <= '0';
      end if;
    end if;
  end process  Energy_Bin_318;   
  
  Energy_Bin_319 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_319   <=  (others =>'0');
		Energy_Bin_Rdy_319 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E319_C1_L and PEAK_C1 <= s_E319_C1_H and Bin_OR = '0') then
         s_Energy_Bin_319 <= s_Energy_Bin_319 +'1';
		 Energy_Bin_Rdy_319 <= '1';
		else
		 s_Energy_Bin_319 <= s_Energy_Bin_319;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_319 <= '0';
      end if;
    end if;
  end process  Energy_Bin_319;       
  
     Energy_Bin_320 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_320   <=  (others =>'0');
		Energy_Bin_Rdy_320 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E320_C1_L and PEAK_C1 <= s_E320_C1_H and Bin_OR = '0') then
         s_Energy_Bin_320 <= s_Energy_Bin_320 +'1';
		 Energy_Bin_Rdy_320 <= '1';
		else
		 s_Energy_Bin_320 <= s_Energy_Bin_320;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_320 <= '0';
      end if;
    end if;
  end process  Energy_Bin_320;    
  
  Energy_Bin_321 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_321   <=  (others =>'0');
		Energy_Bin_Rdy_321 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E321_C1_L and PEAK_C1 <= s_E321_C1_H and Bin_OR = '0') then
         s_Energy_Bin_321 <= s_Energy_Bin_321 +'1';
		 Energy_Bin_Rdy_321 <= '1';
		else
		 s_Energy_Bin_321 <= s_Energy_Bin_321;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_321 <= '0';
      end if;
    end if;
  end process  Energy_Bin_321;   
  
  Energy_Bin_322 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_322   <=  (others =>'0');
	    Energy_Bin_Rdy_322 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E322_C1_L and PEAK_C1 <= s_E322_C1_H and Bin_OR = '0') then
         s_Energy_Bin_322 <= s_Energy_Bin_322 +'1';
		 Energy_Bin_Rdy_322 <= '1';
		else
		 s_Energy_Bin_322 <= s_Energy_Bin_322;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_322 <= '0';
      end if;
    end if;
  end process  Energy_Bin_322;   
  
  Energy_Bin_323 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_323   <=  (others =>'0');
	    Energy_Bin_Rdy_323 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E323_C1_L and PEAK_C1 <= s_E323_C1_H and Bin_OR = '0') then
         s_Energy_Bin_323 <= s_Energy_Bin_323 +'1';
		 Energy_Bin_Rdy_323 <= '1';
		else
		 s_Energy_Bin_323 <= s_Energy_Bin_323;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_323 <= '0';
      end if;
    end if;
  end process  Energy_Bin_323;   
  
  Energy_Bin_324 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_324   <=  (others =>'0');
		Energy_Bin_Rdy_324 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E324_C1_L and PEAK_C1 <= s_E324_C1_H and Bin_OR = '0') then
         s_Energy_Bin_324 <= s_Energy_Bin_324 +'1';
		 Energy_Bin_Rdy_324 <= '1';
		else
		 s_Energy_Bin_324 <= s_Energy_Bin_324;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_324 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_324;   
 
 
  Energy_Bin_325 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_325   <=  (others =>'0');
		Energy_Bin_Rdy_325 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E325_C1_L and PEAK_C1 <= s_E325_C1_H and Bin_OR = '0') then
         s_Energy_Bin_325 <= s_Energy_Bin_325 +'1';
		 Energy_Bin_Rdy_325 <= '1';
		else
		 s_Energy_Bin_325 <= s_Energy_Bin_325;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_325 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_325;  
 
  
  Energy_Bin_326 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_326   <=  (others =>'0');
		Energy_Bin_Rdy_326 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E326_C1_L and PEAK_C1 <= s_E326_C1_H and Bin_OR = '0') then
         s_Energy_Bin_326 <= s_Energy_Bin_326 +'1';
		 Energy_Bin_Rdy_326 <= '1';
		else
		 s_Energy_Bin_326 <= s_Energy_Bin_326;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_326 <= '0';
      end if;
    end if;
  end process  Energy_Bin_326;   
  
 Energy_Bin_327 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_327   <=  (others =>'0');
		Energy_Bin_Rdy_327 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E327_C1_L and PEAK_C1 <= s_E327_C1_H and Bin_OR = '0') then
         s_Energy_Bin_327 <= s_Energy_Bin_327 +'1';
		 Energy_Bin_Rdy_327 <= '1';
		else
		 s_Energy_Bin_327 <= s_Energy_Bin_327;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_327 <= '0';
      end if;
    end if;
  end process  Energy_Bin_327;   
  
  Energy_Bin_328 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_328   <=  (others =>'0');
		Energy_Bin_Rdy_328 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E328_C1_L and PEAK_C1 <= s_E328_C1_H and Bin_OR = '0') then
         s_Energy_Bin_328 <= s_Energy_Bin_328 +'1';
		 Energy_Bin_Rdy_328 <= '1';
		else
		 s_Energy_Bin_328 <= s_Energy_Bin_328;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_328 <= '0';
      end if;
    end if;
  end process  Energy_Bin_328;   
  
  Energy_Bin_329 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_329   <=  (others =>'0');
		Energy_Bin_Rdy_329 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E329_C1_L and PEAK_C1 <= s_E329_C1_H and Bin_OR = '0') then
         s_Energy_Bin_329 <= s_Energy_Bin_329 +'1';
		 Energy_Bin_Rdy_329 <= '1';
		else
		 s_Energy_Bin_329 <= s_Energy_Bin_329;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_329 <= '0';
      end if;
    end if;
  end process  Energy_Bin_329;        
  
     Energy_Bin_330 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_330   <=  (others =>'0');
		Energy_Bin_Rdy_330 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E330_C1_L and PEAK_C1 <= s_E330_C1_H and Bin_OR = '0') then
         s_Energy_Bin_330 <= s_Energy_Bin_330 +'1';
		 Energy_Bin_Rdy_330 <= '1';
		else
		 s_Energy_Bin_330 <= s_Energy_Bin_330;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_330 <= '0';
      end if;
    end if;
  end process  Energy_Bin_330;    
  
  Energy_Bin_331 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_331   <=  (others =>'0');
		Energy_Bin_Rdy_331 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E331_C1_L and PEAK_C1 <= s_E331_C1_H and Bin_OR = '0') then
         s_Energy_Bin_331 <= s_Energy_Bin_331 +'1';
		 Energy_Bin_Rdy_331 <= '1';
		else
		 s_Energy_Bin_331 <= s_Energy_Bin_331;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_331 <= '0';
      end if;
    end if;
  end process  Energy_Bin_331;   
  
  Energy_Bin_332 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_332   <=  (others =>'0');
	    Energy_Bin_Rdy_332 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E332_C1_L and PEAK_C1 <= s_E332_C1_H and Bin_OR = '0') then
         s_Energy_Bin_332 <= s_Energy_Bin_332 +'1';
		 Energy_Bin_Rdy_332 <= '1';
		else
		 s_Energy_Bin_332 <= s_Energy_Bin_332;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_332 <= '0';
      end if;
    end if;
  end process  Energy_Bin_332;   
  
  Energy_Bin_333 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_333   <=  (others =>'0');
	    Energy_Bin_Rdy_333 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E333_C1_L and PEAK_C1 <= s_E333_C1_H and Bin_OR = '0') then
         s_Energy_Bin_333 <= s_Energy_Bin_333 +'1';
		 Energy_Bin_Rdy_333 <= '1';
		else
		 s_Energy_Bin_333 <= s_Energy_Bin_333;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_333 <= '0';
      end if;
    end if;
  end process  Energy_Bin_333;   
  
  Energy_Bin_334 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_334   <=  (others =>'0');
		Energy_Bin_Rdy_334 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E334_C1_L and PEAK_C1 <= s_E334_C1_H and Bin_OR = '0') then
         s_Energy_Bin_334 <= s_Energy_Bin_334 +'1';
		 Energy_Bin_Rdy_334 <= '1';
		else
		 s_Energy_Bin_334 <= s_Energy_Bin_334;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_334 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_334;   
 
 
  Energy_Bin_335 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_335   <=  (others =>'0');
		Energy_Bin_Rdy_335 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E335_C1_L and PEAK_C1 <= s_E335_C1_H and Bin_OR = '0') then
         s_Energy_Bin_335 <= s_Energy_Bin_335 +'1';
		 Energy_Bin_Rdy_335 <= '1';
		else
		 s_Energy_Bin_335 <= s_Energy_Bin_335;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_335 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_335;  
 
  
  Energy_Bin_336 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_336   <=  (others =>'0');
		Energy_Bin_Rdy_336 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E336_C1_L and PEAK_C1 <= s_E336_C1_H and Bin_OR = '0') then
         s_Energy_Bin_336 <= s_Energy_Bin_336 +'1';
		 Energy_Bin_Rdy_336 <= '1';
		else
		 s_Energy_Bin_336 <= s_Energy_Bin_336;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_336 <= '0';
      end if;
    end if;
  end process  Energy_Bin_336;   
  
 Energy_Bin_337 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_337   <=  (others =>'0');
		Energy_Bin_Rdy_337 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E337_C1_L and PEAK_C1 <= s_E337_C1_H and Bin_OR = '0') then
         s_Energy_Bin_337 <= s_Energy_Bin_337 +'1';
		 Energy_Bin_Rdy_337 <= '1';
		else
		 s_Energy_Bin_337 <= s_Energy_Bin_337;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_337 <= '0';
      end if;
    end if;
  end process  Energy_Bin_337;   
  
  Energy_Bin_338 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_338   <=  (others =>'0');
		Energy_Bin_Rdy_338 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E338_C1_L and PEAK_C1 <= s_E338_C1_H and Bin_OR = '0') then
         s_Energy_Bin_338 <= s_Energy_Bin_338 +'1';
		 Energy_Bin_Rdy_338 <= '1';
		else
		 s_Energy_Bin_338 <= s_Energy_Bin_338;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_338 <= '0';
      end if;
    end if;
  end process  Energy_Bin_338;   
  
  Energy_Bin_339 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_339   <=  (others =>'0');
		Energy_Bin_Rdy_339 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E339_C1_L and PEAK_C1 <= s_E339_C1_H and Bin_OR = '0') then
         s_Energy_Bin_339 <= s_Energy_Bin_339 +'1';
		 Energy_Bin_Rdy_339 <= '1';
		else
		 s_Energy_Bin_339 <= s_Energy_Bin_339;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_339 <= '0';
      end if;
    end if;
  end process  Energy_Bin_339;         
  
     Energy_Bin_340 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_340   <=  (others =>'0');
		Energy_Bin_Rdy_340 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E340_C1_L and PEAK_C1 <= s_E340_C1_H and Bin_OR = '0') then
         s_Energy_Bin_340 <= s_Energy_Bin_340 +'1';
		 Energy_Bin_Rdy_340 <= '1';
		else
		 s_Energy_Bin_340 <= s_Energy_Bin_340;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_340 <= '0';
      end if;
    end if;
  end process  Energy_Bin_340;    
  
  Energy_Bin_341 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_341   <=  (others =>'0');
		Energy_Bin_Rdy_341 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E341_C1_L and PEAK_C1 <= s_E341_C1_H and Bin_OR = '0') then
         s_Energy_Bin_341 <= s_Energy_Bin_341 +'1';
		 Energy_Bin_Rdy_341 <= '1';
		else
		 s_Energy_Bin_341 <= s_Energy_Bin_341;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_341 <= '0';
      end if;
    end if;
  end process  Energy_Bin_341;   
  
  Energy_Bin_342 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_342   <=  (others =>'0');
	    Energy_Bin_Rdy_342 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E342_C1_L and PEAK_C1 <= s_E342_C1_H and Bin_OR = '0') then
         s_Energy_Bin_342 <= s_Energy_Bin_342 +'1';
		 Energy_Bin_Rdy_342 <= '1';
		else
		 s_Energy_Bin_342 <= s_Energy_Bin_342;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_342 <= '0';
      end if;
    end if;
  end process  Energy_Bin_342;   
  
  Energy_Bin_343 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_343   <=  (others =>'0');
	    Energy_Bin_Rdy_343 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E343_C1_L and PEAK_C1 <= s_E343_C1_H and Bin_OR = '0') then
         s_Energy_Bin_343 <= s_Energy_Bin_343 +'1';
		 Energy_Bin_Rdy_343 <= '1';
		else
		 s_Energy_Bin_343 <= s_Energy_Bin_343;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_343 <= '0';
      end if;
    end if;
  end process  Energy_Bin_343;   
  
  Energy_Bin_344 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_344   <=  (others =>'0');
		Energy_Bin_Rdy_344 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E344_C1_L and PEAK_C1 <= s_E344_C1_H and Bin_OR = '0') then
         s_Energy_Bin_344 <= s_Energy_Bin_344 +'1';
		 Energy_Bin_Rdy_344 <= '1';
		else
		 s_Energy_Bin_344 <= s_Energy_Bin_344;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_344 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_344;   
 
 
  Energy_Bin_345 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_345   <=  (others =>'0');
		Energy_Bin_Rdy_345 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E345_C1_L and PEAK_C1 <= s_E345_C1_H and Bin_OR = '0') then
         s_Energy_Bin_345 <= s_Energy_Bin_345 +'1';
		 Energy_Bin_Rdy_345 <= '1';
		else
		 s_Energy_Bin_345 <= s_Energy_Bin_345;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_345 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_345;  
 
  
  Energy_Bin_346 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_346   <=  (others =>'0');
		Energy_Bin_Rdy_346 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E346_C1_L and PEAK_C1 <= s_E346_C1_H and Bin_OR = '0') then
         s_Energy_Bin_346 <= s_Energy_Bin_346 +'1';
		 Energy_Bin_Rdy_346 <= '1';
		else
		 s_Energy_Bin_346 <= s_Energy_Bin_346;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_346 <= '0';
      end if;
    end if;
  end process  Energy_Bin_346;   
  
 Energy_Bin_347 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_347   <=  (others =>'0');
		Energy_Bin_Rdy_347 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E347_C1_L and PEAK_C1 <= s_E347_C1_H and Bin_OR = '0') then
         s_Energy_Bin_347 <= s_Energy_Bin_347 +'1';
		 Energy_Bin_Rdy_347 <= '1';
		else
		 s_Energy_Bin_347 <= s_Energy_Bin_347;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_347 <= '0';
      end if;
    end if;
  end process  Energy_Bin_347;   
  
  Energy_Bin_348 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_348   <=  (others =>'0');
		Energy_Bin_Rdy_348 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E348_C1_L and PEAK_C1 <= s_E348_C1_H and Bin_OR = '0') then
         s_Energy_Bin_348 <= s_Energy_Bin_348 +'1';
		 Energy_Bin_Rdy_348 <= '1';
		else
		 s_Energy_Bin_348 <= s_Energy_Bin_348;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_348 <= '0';
      end if;
    end if;
  end process  Energy_Bin_348;   
  
  Energy_Bin_349 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_349   <=  (others =>'0');
		Energy_Bin_Rdy_349 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E349_C1_L and PEAK_C1 <= s_E349_C1_H and Bin_OR = '0') then
         s_Energy_Bin_349 <= s_Energy_Bin_349 +'1';
		 Energy_Bin_Rdy_349 <= '1';
		else
		 s_Energy_Bin_349 <= s_Energy_Bin_349;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_349 <= '0';
      end if;
    end if;
  end process  Energy_Bin_349;          
  
  
     Energy_Bin_350 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_350   <=  (others =>'0');
		Energy_Bin_Rdy_350 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E350_C1_L and PEAK_C1 <= s_E350_C1_H and Bin_OR = '0') then
         s_Energy_Bin_350 <= s_Energy_Bin_350 +'1';
		 Energy_Bin_Rdy_350 <= '1';
		else
		 s_Energy_Bin_350 <= s_Energy_Bin_350;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_350 <= '0';
      end if;
    end if;
  end process  Energy_Bin_350;    
  
  Energy_Bin_351 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_351   <=  (others =>'0');
		Energy_Bin_Rdy_351 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E351_C1_L and PEAK_C1 <= s_E351_C1_H and Bin_OR = '0') then
         s_Energy_Bin_351 <= s_Energy_Bin_351 +'1';
		 Energy_Bin_Rdy_351 <= '1';
		else
		 s_Energy_Bin_351 <= s_Energy_Bin_351;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_351 <= '0';
      end if;
    end if;
  end process  Energy_Bin_351;   
  
  Energy_Bin_352 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_352   <=  (others =>'0');
	    Energy_Bin_Rdy_352 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E352_C1_L and PEAK_C1 <= s_E352_C1_H and Bin_OR = '0') then
         s_Energy_Bin_352 <= s_Energy_Bin_352 +'1';
		 Energy_Bin_Rdy_352 <= '1';
		else
		 s_Energy_Bin_352 <= s_Energy_Bin_352;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_352 <= '0';
      end if;
    end if;
  end process  Energy_Bin_352;   
  
  Energy_Bin_353 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_353   <=  (others =>'0');
	    Energy_Bin_Rdy_353 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E353_C1_L and PEAK_C1 <= s_E353_C1_H and Bin_OR = '0') then
         s_Energy_Bin_353 <= s_Energy_Bin_353 +'1';
		 Energy_Bin_Rdy_353 <= '1';
		else
		 s_Energy_Bin_353 <= s_Energy_Bin_353;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_353 <= '0';
      end if;
    end if;
  end process  Energy_Bin_353;   
  
  Energy_Bin_354 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_354   <=  (others =>'0');
		Energy_Bin_Rdy_354 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E354_C1_L and PEAK_C1 <= s_E354_C1_H and Bin_OR = '0') then
         s_Energy_Bin_354 <= s_Energy_Bin_354 +'1';
		 Energy_Bin_Rdy_354 <= '1';
		else
		 s_Energy_Bin_354 <= s_Energy_Bin_354;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_354 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_354;   
 
 
  Energy_Bin_355 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_355   <=  (others =>'0');
		Energy_Bin_Rdy_355 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E355_C1_L and PEAK_C1 <= s_E355_C1_H and Bin_OR = '0') then
         s_Energy_Bin_355 <= s_Energy_Bin_355 +'1';
		 Energy_Bin_Rdy_355 <= '1';
		else
		 s_Energy_Bin_355 <= s_Energy_Bin_355;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_355 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_355;  
 
  
  Energy_Bin_356 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_356   <=  (others =>'0');
		Energy_Bin_Rdy_356 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E356_C1_L and PEAK_C1 <= s_E356_C1_H and Bin_OR = '0') then
         s_Energy_Bin_356 <= s_Energy_Bin_356 +'1';
		 Energy_Bin_Rdy_356 <= '1';
		else
		 s_Energy_Bin_356 <= s_Energy_Bin_356;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_356 <= '0';
      end if;
    end if;
  end process  Energy_Bin_356;   
  
 Energy_Bin_357 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_357   <=  (others =>'0');
		Energy_Bin_Rdy_357 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E357_C1_L and PEAK_C1 <= s_E357_C1_H and Bin_OR = '0') then
         s_Energy_Bin_357 <= s_Energy_Bin_357 +'1';
		 Energy_Bin_Rdy_357 <= '1';
		else
		 s_Energy_Bin_357 <= s_Energy_Bin_357;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_357 <= '0';
      end if;
    end if;
  end process  Energy_Bin_357;   
  
  Energy_Bin_358 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_358   <=  (others =>'0');
		Energy_Bin_Rdy_358 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E358_C1_L and PEAK_C1 <= s_E358_C1_H and Bin_OR = '0') then
         s_Energy_Bin_358 <= s_Energy_Bin_358 +'1';
		 Energy_Bin_Rdy_358 <= '1';
		else
		 s_Energy_Bin_358 <= s_Energy_Bin_358;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_358 <= '0';
      end if;
    end if;
  end process  Energy_Bin_358;   
  
  Energy_Bin_359 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_359   <=  (others =>'0');
		Energy_Bin_Rdy_359 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E359_C1_L and PEAK_C1 <= s_E359_C1_H and Bin_OR = '0') then
         s_Energy_Bin_359 <= s_Energy_Bin_359 +'1';
		 Energy_Bin_Rdy_359 <= '1';
		else
		 s_Energy_Bin_359 <= s_Energy_Bin_359;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_359 <= '0';
      end if;
    end if;
  end process  Energy_Bin_359;           
  
     Energy_Bin_360 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_360   <=  (others =>'0');
		Energy_Bin_Rdy_360 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E360_C1_L and PEAK_C1 <= s_E360_C1_H and Bin_OR = '0') then
         s_Energy_Bin_360 <= s_Energy_Bin_360 +'1';
		 Energy_Bin_Rdy_360 <= '1';
		else
		 s_Energy_Bin_360 <= s_Energy_Bin_360;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_360 <= '0';
      end if;
    end if;
  end process  Energy_Bin_360;    
  
  Energy_Bin_361 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_361   <=  (others =>'0');
		Energy_Bin_Rdy_361 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E361_C1_L and PEAK_C1 <= s_E361_C1_H and Bin_OR = '0') then
         s_Energy_Bin_361 <= s_Energy_Bin_361 +'1';
		 Energy_Bin_Rdy_361 <= '1';
		else
		 s_Energy_Bin_361 <= s_Energy_Bin_361;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_361 <= '0';
      end if;
    end if;
  end process  Energy_Bin_361;   
  
  Energy_Bin_362 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_362   <=  (others =>'0');
	    Energy_Bin_Rdy_362 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E362_C1_L and PEAK_C1 <= s_E362_C1_H and Bin_OR = '0') then
         s_Energy_Bin_362 <= s_Energy_Bin_362 +'1';
		 Energy_Bin_Rdy_362 <= '1';
		else
		 s_Energy_Bin_362 <= s_Energy_Bin_362;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_362 <= '0';
      end if;
    end if;
  end process  Energy_Bin_362;   
  
  Energy_Bin_363 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_363   <=  (others =>'0');
	    Energy_Bin_Rdy_363 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E363_C1_L and PEAK_C1 <= s_E363_C1_H and Bin_OR = '0') then
         s_Energy_Bin_363 <= s_Energy_Bin_363 +'1';
		 Energy_Bin_Rdy_363 <= '1';
		else
		 s_Energy_Bin_363 <= s_Energy_Bin_363;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_363 <= '0';
      end if;
    end if;
  end process  Energy_Bin_363;   
  
  Energy_Bin_364 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_364   <=  (others =>'0');
		Energy_Bin_Rdy_364 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E364_C1_L and PEAK_C1 <= s_E364_C1_H and Bin_OR = '0') then
         s_Energy_Bin_364 <= s_Energy_Bin_364 +'1';
		 Energy_Bin_Rdy_364 <= '1';
		else
		 s_Energy_Bin_364 <= s_Energy_Bin_364;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_364 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_364;   
 
 
  Energy_Bin_365 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_365   <=  (others =>'0');
		Energy_Bin_Rdy_365 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E365_C1_L and PEAK_C1 <= s_E365_C1_H and Bin_OR = '0') then
         s_Energy_Bin_365 <= s_Energy_Bin_365 +'1';
		 Energy_Bin_Rdy_365 <= '1';
		else
		 s_Energy_Bin_365 <= s_Energy_Bin_365;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_365 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_365;  
 
  
  Energy_Bin_366 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_366   <=  (others =>'0');
		Energy_Bin_Rdy_366 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E366_C1_L and PEAK_C1 <= s_E366_C1_H and Bin_OR = '0') then
         s_Energy_Bin_366 <= s_Energy_Bin_366 +'1';
		 Energy_Bin_Rdy_366 <= '1';
		else
		 s_Energy_Bin_366 <= s_Energy_Bin_366;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_366 <= '0';
      end if;
    end if;
  end process  Energy_Bin_366;   
  
 Energy_Bin_367 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_367   <=  (others =>'0');
		Energy_Bin_Rdy_367 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E367_C1_L and PEAK_C1 <= s_E367_C1_H and Bin_OR = '0') then
         s_Energy_Bin_367 <= s_Energy_Bin_367 +'1';
		 Energy_Bin_Rdy_367 <= '1';
		else
		 s_Energy_Bin_367 <= s_Energy_Bin_367;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_367 <= '0';
      end if;
    end if;
  end process  Energy_Bin_367;   
  
  Energy_Bin_368 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_368   <=  (others =>'0');
		Energy_Bin_Rdy_368 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E368_C1_L and PEAK_C1 <= s_E368_C1_H and Bin_OR = '0') then
         s_Energy_Bin_368 <= s_Energy_Bin_368 +'1';
		 Energy_Bin_Rdy_368 <= '1';
		else
		 s_Energy_Bin_368 <= s_Energy_Bin_368;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_368 <= '0';
      end if;
    end if;
  end process  Energy_Bin_368;   
  
  Energy_Bin_369 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_369   <=  (others =>'0');
		Energy_Bin_Rdy_369 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E369_C1_L and PEAK_C1 <= s_E369_C1_H and Bin_OR = '0') then
         s_Energy_Bin_369 <= s_Energy_Bin_369 +'1';
		 Energy_Bin_Rdy_369 <= '1';
		else
		 s_Energy_Bin_369 <= s_Energy_Bin_369;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_369 <= '0';
      end if;
    end if;
  end process  Energy_Bin_369;         
  
     Energy_Bin_370 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_370   <=  (others =>'0');
		Energy_Bin_Rdy_370 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E370_C1_L and PEAK_C1 <= s_E370_C1_H and Bin_OR = '0') then
         s_Energy_Bin_370 <= s_Energy_Bin_370 +'1';
		 Energy_Bin_Rdy_370 <= '1';
		else
		 s_Energy_Bin_370 <= s_Energy_Bin_370;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_370 <= '0';
      end if;
    end if;
  end process  Energy_Bin_370;    
  
  Energy_Bin_371 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_371   <=  (others =>'0');
		Energy_Bin_Rdy_371 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E371_C1_L and PEAK_C1 <= s_E371_C1_H and Bin_OR = '0') then
         s_Energy_Bin_371 <= s_Energy_Bin_371 +'1';
		 Energy_Bin_Rdy_371 <= '1';
		else
		 s_Energy_Bin_371 <= s_Energy_Bin_371;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_371 <= '0';
      end if;
    end if;
  end process  Energy_Bin_371;   
  
  Energy_Bin_372 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_372   <=  (others =>'0');
	    Energy_Bin_Rdy_372 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E372_C1_L and PEAK_C1 <= s_E372_C1_H and Bin_OR = '0') then
         s_Energy_Bin_372 <= s_Energy_Bin_372 +'1';
		 Energy_Bin_Rdy_372 <= '1';
		else
		 s_Energy_Bin_372 <= s_Energy_Bin_372;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_372 <= '0';
      end if;
    end if;
  end process  Energy_Bin_372;   
  
  Energy_Bin_373 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_373   <=  (others =>'0');
	    Energy_Bin_Rdy_373 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E373_C1_L and PEAK_C1 <= s_E373_C1_H and Bin_OR = '0') then
         s_Energy_Bin_373 <= s_Energy_Bin_373 +'1';
		 Energy_Bin_Rdy_373 <= '1';
		else
		 s_Energy_Bin_373 <= s_Energy_Bin_373;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_373 <= '0';
      end if;
    end if;
  end process  Energy_Bin_373;   
  
  Energy_Bin_374 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_374   <=  (others =>'0');
		Energy_Bin_Rdy_374 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E374_C1_L and PEAK_C1 <= s_E374_C1_H and Bin_OR = '0') then
         s_Energy_Bin_374 <= s_Energy_Bin_374 +'1';
		 Energy_Bin_Rdy_374 <= '1';
		else
		 s_Energy_Bin_374 <= s_Energy_Bin_374;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_374 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_374;   
 
 
  Energy_Bin_375 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_375   <=  (others =>'0');
		Energy_Bin_Rdy_375 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E375_C1_L and PEAK_C1 <= s_E375_C1_H and Bin_OR = '0') then
         s_Energy_Bin_375 <= s_Energy_Bin_375 +'1';
		 Energy_Bin_Rdy_375 <= '1';
		else
		 s_Energy_Bin_375 <= s_Energy_Bin_375;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_375 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_375;  
 
  
  Energy_Bin_376 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_376   <=  (others =>'0');
		Energy_Bin_Rdy_376 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E376_C1_L and PEAK_C1 <= s_E376_C1_H and Bin_OR = '0') then
         s_Energy_Bin_376 <= s_Energy_Bin_376 +'1';
		 Energy_Bin_Rdy_376 <= '1';
		else
		 s_Energy_Bin_376 <= s_Energy_Bin_376;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_376 <= '0';
      end if;
    end if;
  end process  Energy_Bin_376;   
  
 Energy_Bin_377 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_377   <=  (others =>'0');
		Energy_Bin_Rdy_377 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E377_C1_L and PEAK_C1 <= s_E377_C1_H and Bin_OR = '0') then
         s_Energy_Bin_377 <= s_Energy_Bin_377 +'1';
		 Energy_Bin_Rdy_377 <= '1';
		else
		 s_Energy_Bin_377 <= s_Energy_Bin_377;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_377 <= '0';
      end if;
    end if;
  end process  Energy_Bin_377;   
  
  Energy_Bin_378 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_378   <=  (others =>'0');
		Energy_Bin_Rdy_378 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E378_C1_L and PEAK_C1 <= s_E378_C1_H and Bin_OR = '0') then
         s_Energy_Bin_378 <= s_Energy_Bin_378 +'1';
		 Energy_Bin_Rdy_378 <= '1';
		else
		 s_Energy_Bin_378 <= s_Energy_Bin_378;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_378 <= '0';
      end if;
    end if;
  end process  Energy_Bin_378;   
  
  Energy_Bin_379 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_379   <=  (others =>'0');
		Energy_Bin_Rdy_379 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E379_C1_L and PEAK_C1 <= s_E379_C1_H and Bin_OR = '0') then
         s_Energy_Bin_379 <= s_Energy_Bin_379 +'1';
		 Energy_Bin_Rdy_379 <= '1';
		else
		 s_Energy_Bin_379 <= s_Energy_Bin_379;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_379 <= '0';
      end if;
    end if;
  end process  Energy_Bin_379;       
  
     Energy_Bin_380 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_380   <=  (others =>'0');
		Energy_Bin_Rdy_380 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E380_C1_L and PEAK_C1 <= s_E380_C1_H and Bin_OR = '0') then
         s_Energy_Bin_380 <= s_Energy_Bin_380 +'1';
		 Energy_Bin_Rdy_380 <= '1';
		else
		 s_Energy_Bin_380 <= s_Energy_Bin_380;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_380 <= '0';
      end if;
    end if;
  end process  Energy_Bin_380;    
  
  Energy_Bin_381 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_381   <=  (others =>'0');
		Energy_Bin_Rdy_381 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E381_C1_L and PEAK_C1 <= s_E381_C1_H and Bin_OR = '0') then
         s_Energy_Bin_381 <= s_Energy_Bin_381 +'1';
		 Energy_Bin_Rdy_381 <= '1';
		else
		 s_Energy_Bin_381 <= s_Energy_Bin_381;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_381 <= '0';
      end if;
    end if;
  end process  Energy_Bin_381;   
  
  Energy_Bin_382 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_382   <=  (others =>'0');
	    Energy_Bin_Rdy_382 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E382_C1_L and PEAK_C1 <= s_E382_C1_H and Bin_OR = '0') then
         s_Energy_Bin_382 <= s_Energy_Bin_382 +'1';
		 Energy_Bin_Rdy_382 <= '1';
		else
		 s_Energy_Bin_382 <= s_Energy_Bin_382;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_382 <= '0';
      end if;
    end if;
  end process  Energy_Bin_382;   
  
  Energy_Bin_383 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_383   <=  (others =>'0');
	    Energy_Bin_Rdy_383 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E383_C1_L and PEAK_C1 <= s_E383_C1_H and Bin_OR = '0') then
         s_Energy_Bin_383 <= s_Energy_Bin_383 +'1';
		 Energy_Bin_Rdy_383 <= '1';
		else
		 s_Energy_Bin_383 <= s_Energy_Bin_383;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_383 <= '0';
      end if;
    end if;
  end process  Energy_Bin_383;   
  
  Energy_Bin_384 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_384   <=  (others =>'0');
		Energy_Bin_Rdy_384 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E384_C1_L and PEAK_C1 <= s_E384_C1_H and Bin_OR = '0') then
         s_Energy_Bin_384 <= s_Energy_Bin_384 +'1';
		 Energy_Bin_Rdy_384 <= '1';
		else
		 s_Energy_Bin_384 <= s_Energy_Bin_384;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_384 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_384;   
 
 
  Energy_Bin_385 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_385   <=  (others =>'0');
		Energy_Bin_Rdy_385 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E385_C1_L and PEAK_C1 <= s_E385_C1_H and Bin_OR = '0') then
         s_Energy_Bin_385 <= s_Energy_Bin_385 +'1';
		 Energy_Bin_Rdy_385 <= '1';
		else
		 s_Energy_Bin_385 <= s_Energy_Bin_385;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_385 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_385;  
 
  
  Energy_Bin_386 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_386   <=  (others =>'0');
		Energy_Bin_Rdy_386 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E386_C1_L and PEAK_C1 <= s_E386_C1_H and Bin_OR = '0') then
         s_Energy_Bin_386 <= s_Energy_Bin_386 +'1';
		 Energy_Bin_Rdy_386 <= '1';
		else
		 s_Energy_Bin_386 <= s_Energy_Bin_386;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_386 <= '0';
      end if;
    end if;
  end process  Energy_Bin_386;   
  
 Energy_Bin_387 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_387   <=  (others =>'0');
		Energy_Bin_Rdy_387 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E387_C1_L and PEAK_C1 <= s_E387_C1_H and Bin_OR = '0') then
         s_Energy_Bin_387 <= s_Energy_Bin_387 +'1';
		 Energy_Bin_Rdy_387 <= '1';
		else
		 s_Energy_Bin_387 <= s_Energy_Bin_387;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_387 <= '0';
      end if;
    end if;
  end process  Energy_Bin_387;   
  
  Energy_Bin_388 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_388   <=  (others =>'0');
		Energy_Bin_Rdy_388 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E388_C1_L and PEAK_C1 <= s_E388_C1_H and Bin_OR = '0') then
         s_Energy_Bin_388 <= s_Energy_Bin_388 +'1';
		 Energy_Bin_Rdy_388 <= '1';
		else
		 s_Energy_Bin_388 <= s_Energy_Bin_388;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_388 <= '0';
      end if;
    end if;
  end process  Energy_Bin_388;   
  
  Energy_Bin_389 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_389   <=  (others =>'0');
		Energy_Bin_Rdy_389 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E389_C1_L and PEAK_C1 <= s_E389_C1_H and Bin_OR = '0') then
         s_Energy_Bin_389 <= s_Energy_Bin_389 +'1';
		 Energy_Bin_Rdy_389 <= '1';
		else
		 s_Energy_Bin_389 <= s_Energy_Bin_389;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_389 <= '0';
      end if;
    end if;
  end process  Energy_Bin_389;      
  
     Energy_Bin_390 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_390   <=  (others =>'0');
		Energy_Bin_Rdy_390 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E390_C1_L and PEAK_C1 <= s_E390_C1_H and Bin_OR = '0') then
         s_Energy_Bin_390 <= s_Energy_Bin_390 +'1';
		 Energy_Bin_Rdy_390 <= '1';
		else
		 s_Energy_Bin_390 <= s_Energy_Bin_390;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_390 <= '0';
      end if;
    end if;
  end process  Energy_Bin_390;    
  
  Energy_Bin_391 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_391   <=  (others =>'0');
		Energy_Bin_Rdy_391 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E391_C1_L and PEAK_C1 <= s_E391_C1_H and Bin_OR = '0') then
         s_Energy_Bin_391 <= s_Energy_Bin_391 +'1';
		 Energy_Bin_Rdy_391 <= '1';
		else
		 s_Energy_Bin_391 <= s_Energy_Bin_391;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_391 <= '0';
      end if;
    end if;
  end process  Energy_Bin_391;   
  
  Energy_Bin_392 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_392   <=  (others =>'0');
	    Energy_Bin_Rdy_392 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E392_C1_L and PEAK_C1 <= s_E392_C1_H and Bin_OR = '0') then
         s_Energy_Bin_392 <= s_Energy_Bin_392 +'1';
		 Energy_Bin_Rdy_392 <= '1';
		else
		 s_Energy_Bin_392 <= s_Energy_Bin_392;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_392 <= '0';
      end if;
    end if;
  end process  Energy_Bin_392;   
  
  Energy_Bin_393 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_393   <=  (others =>'0');
	    Energy_Bin_Rdy_393 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E393_C1_L and PEAK_C1 <= s_E393_C1_H and Bin_OR = '0') then
         s_Energy_Bin_393 <= s_Energy_Bin_393 +'1';
		 Energy_Bin_Rdy_393 <= '1';
		else
		 s_Energy_Bin_393 <= s_Energy_Bin_393;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_393 <= '0';
      end if;
    end if;
  end process  Energy_Bin_393;   
  
  Energy_Bin_394 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_394   <=  (others =>'0');
		Energy_Bin_Rdy_394 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E394_C1_L and PEAK_C1 <= s_E394_C1_H and Bin_OR = '0') then
         s_Energy_Bin_394 <= s_Energy_Bin_394 +'1';
		 Energy_Bin_Rdy_394 <= '1';
		else
		 s_Energy_Bin_394 <= s_Energy_Bin_394;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_394 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_394;   
 
 
  Energy_Bin_395 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_395   <=  (others =>'0');
		Energy_Bin_Rdy_395 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E395_C1_L and PEAK_C1 <= s_E395_C1_H and Bin_OR = '0') then
         s_Energy_Bin_395 <= s_Energy_Bin_395 +'1';
		 Energy_Bin_Rdy_395 <= '1';
		else
		 s_Energy_Bin_395 <= s_Energy_Bin_395;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_395 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_395;  
 
  
  Energy_Bin_396 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_396   <=  (others =>'0');
		Energy_Bin_Rdy_396 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E396_C1_L and PEAK_C1 <= s_E396_C1_H and Bin_OR = '0') then
         s_Energy_Bin_396 <= s_Energy_Bin_396 +'1';
		 Energy_Bin_Rdy_396 <= '1';
		else
		 s_Energy_Bin_396 <= s_Energy_Bin_396;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_396 <= '0';
      end if;
    end if;
  end process  Energy_Bin_396;   
  
 Energy_Bin_397 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_397   <=  (others =>'0');
		Energy_Bin_Rdy_397 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E397_C1_L and PEAK_C1 <= s_E397_C1_H and Bin_OR = '0') then
         s_Energy_Bin_397 <= s_Energy_Bin_397 +'1';
		 Energy_Bin_Rdy_397 <= '1';
		else
		 s_Energy_Bin_397 <= s_Energy_Bin_397;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_397 <= '0';
      end if;
    end if;
  end process  Energy_Bin_397;   
  
  Energy_Bin_398 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_398   <=  (others =>'0');
		Energy_Bin_Rdy_398 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E398_C1_L and PEAK_C1 <= s_E398_C1_H and Bin_OR = '0') then
         s_Energy_Bin_398 <= s_Energy_Bin_398 +'1';
		 Energy_Bin_Rdy_398 <= '1';
		else
		 s_Energy_Bin_398 <= s_Energy_Bin_398;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_398 <= '0';
      end if;
    end if;
  end process  Energy_Bin_398;   
  
  Energy_Bin_399 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_399   <=  (others =>'0');
		Energy_Bin_Rdy_399 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E399_C1_L and PEAK_C1 <= s_E399_C1_H and Bin_OR = '0') then
         s_Energy_Bin_399 <= s_Energy_Bin_399 +'1';
		 Energy_Bin_Rdy_399 <= '1';
		else
		 s_Energy_Bin_399 <= s_Energy_Bin_399;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_399 <= '0';
      end if;
    end if;
  end process  Energy_Bin_399;      

    Energy_Bin_400 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_400   <=  (others =>'0');
		Energy_Bin_Rdy_400 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E400_C1_L and PEAK_C1 <= s_E400_C1_H and Bin_OR = '0') then
         s_Energy_Bin_400 <= s_Energy_Bin_400 +'1';
		 Energy_Bin_Rdy_400 <= '1';
		else
		 s_Energy_Bin_400 <= s_Energy_Bin_400;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_400 <= '0';
      end if;
    end if;
  end process  Energy_Bin_400;    
  
  Energy_Bin_401 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_401   <=  (others =>'0');
		Energy_Bin_Rdy_401 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E401_C1_L and PEAK_C1 <= s_E401_C1_H and Bin_OR = '0') then
         s_Energy_Bin_401 <= s_Energy_Bin_401 +'1';
		 Energy_Bin_Rdy_401 <= '1';
		else
		 s_Energy_Bin_401 <= s_Energy_Bin_401;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_401 <= '0';
      end if;
    end if;
  end process  Energy_Bin_401;   
  
  Energy_Bin_402 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_402   <=  (others =>'0');
	    Energy_Bin_Rdy_402 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E402_C1_L and PEAK_C1 <= s_E402_C1_H and Bin_OR = '0') then
         s_Energy_Bin_402 <= s_Energy_Bin_402 +'1';
		 Energy_Bin_Rdy_402 <= '1';
		else
		 s_Energy_Bin_402 <= s_Energy_Bin_402;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_402 <= '0';
      end if;
    end if;
  end process  Energy_Bin_402;   
  
  Energy_Bin_403 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_403   <=  (others =>'0');
	    Energy_Bin_Rdy_403 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E403_C1_L and PEAK_C1 <= s_E403_C1_H and Bin_OR = '0') then
         s_Energy_Bin_403 <= s_Energy_Bin_403 +'1';
		 Energy_Bin_Rdy_403 <= '1';
		else
		 s_Energy_Bin_403 <= s_Energy_Bin_403;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_403 <= '0';
      end if;
    end if;
  end process  Energy_Bin_403;   
  
  Energy_Bin_404 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_404   <=  (others =>'0');
		Energy_Bin_Rdy_404 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E404_C1_L and PEAK_C1 <= s_E404_C1_H and Bin_OR = '0') then
         s_Energy_Bin_404 <= s_Energy_Bin_404 +'1';
		 Energy_Bin_Rdy_404 <= '1';
		else
		 s_Energy_Bin_404 <= s_Energy_Bin_404;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_404 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_404;   
 
 
  Energy_Bin_405 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_405   <=  (others =>'0');
		Energy_Bin_Rdy_405 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E405_C1_L and PEAK_C1 <= s_E405_C1_H and Bin_OR = '0') then
         s_Energy_Bin_405 <= s_Energy_Bin_405 +'1';
		 Energy_Bin_Rdy_405 <= '1';
		else
		 s_Energy_Bin_405 <= s_Energy_Bin_405;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_405 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_405;  
 
  
  Energy_Bin_406 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_406   <=  (others =>'0');
		Energy_Bin_Rdy_406 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E406_C1_L and PEAK_C1 <= s_E406_C1_H and Bin_OR = '0') then
         s_Energy_Bin_406 <= s_Energy_Bin_406 +'1';
		 Energy_Bin_Rdy_406 <= '1';
		else
		 s_Energy_Bin_406 <= s_Energy_Bin_406;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_406 <= '0';
      end if;
    end if;
  end process  Energy_Bin_406;   
  
 Energy_Bin_407 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_407   <=  (others =>'0');
		Energy_Bin_Rdy_407 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E407_C1_L and PEAK_C1 <= s_E407_C1_H and Bin_OR = '0') then
         s_Energy_Bin_407 <= s_Energy_Bin_407 +'1';
		 Energy_Bin_Rdy_407 <= '1';
		else
		 s_Energy_Bin_407 <= s_Energy_Bin_407;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_407 <= '0';
      end if;
    end if;
  end process  Energy_Bin_407;   
  
  Energy_Bin_408 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_408   <=  (others =>'0');
		Energy_Bin_Rdy_408 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E408_C1_L and PEAK_C1 <= s_E408_C1_H and Bin_OR = '0') then
         s_Energy_Bin_408 <= s_Energy_Bin_408 +'1';
		 Energy_Bin_Rdy_408 <= '1';
		else
		 s_Energy_Bin_408 <= s_Energy_Bin_408;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_408 <= '0';
      end if;
    end if;
  end process  Energy_Bin_408;   
  
  Energy_Bin_409 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_409   <=  (others =>'0');
		Energy_Bin_Rdy_409 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E409_C1_L and PEAK_C1 <= s_E409_C1_H and Bin_OR = '0') then
         s_Energy_Bin_409 <= s_Energy_Bin_409 +'1';
		 Energy_Bin_Rdy_409 <= '1';
		else
		 s_Energy_Bin_409 <= s_Energy_Bin_409;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_409 <= '0';
      end if;
    end if;
  end process  Energy_Bin_409;      
  
     Energy_Bin_410 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_410   <=  (others =>'0');
		Energy_Bin_Rdy_410 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E410_C1_L and PEAK_C1 <= s_E410_C1_H and Bin_OR = '0') then
         s_Energy_Bin_410 <= s_Energy_Bin_410 +'1';
		 Energy_Bin_Rdy_410 <= '1';
		else
		 s_Energy_Bin_410 <= s_Energy_Bin_410;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_410 <= '0';
      end if;
    end if;
  end process  Energy_Bin_410;    
  
  Energy_Bin_411 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_411   <=  (others =>'0');
		Energy_Bin_Rdy_411 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E411_C1_L and PEAK_C1 <= s_E411_C1_H and Bin_OR = '0') then
         s_Energy_Bin_411 <= s_Energy_Bin_411 +'1';
		 Energy_Bin_Rdy_411 <= '1';
		else
		 s_Energy_Bin_411 <= s_Energy_Bin_411;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_411 <= '0';
      end if;
    end if;
  end process  Energy_Bin_411;   
  
  Energy_Bin_412 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_412   <=  (others =>'0');
	    Energy_Bin_Rdy_412 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E412_C1_L and PEAK_C1 <= s_E412_C1_H and Bin_OR = '0') then
         s_Energy_Bin_412 <= s_Energy_Bin_412 +'1';
		 Energy_Bin_Rdy_412 <= '1';
		else
		 s_Energy_Bin_412 <= s_Energy_Bin_412;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_412 <= '0';
      end if;
    end if;
  end process  Energy_Bin_412;   
  
  Energy_Bin_413 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_413   <=  (others =>'0');
	    Energy_Bin_Rdy_413 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E413_C1_L and PEAK_C1 <= s_E413_C1_H and Bin_OR = '0') then
         s_Energy_Bin_413 <= s_Energy_Bin_413 +'1';
		 Energy_Bin_Rdy_413 <= '1';
		else
		 s_Energy_Bin_413 <= s_Energy_Bin_413;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_413 <= '0';
      end if;
    end if;
  end process  Energy_Bin_413;   
  
  Energy_Bin_414 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_414   <=  (others =>'0');
		Energy_Bin_Rdy_414 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E414_C1_L and PEAK_C1 <= s_E414_C1_H and Bin_OR = '0') then
         s_Energy_Bin_414 <= s_Energy_Bin_414 +'1';
		 Energy_Bin_Rdy_414 <= '1';
		else
		 s_Energy_Bin_414 <= s_Energy_Bin_414;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_414 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_414;   
 
 
  Energy_Bin_415 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_415   <=  (others =>'0');
		Energy_Bin_Rdy_415 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E415_C1_L and PEAK_C1 <= s_E415_C1_H and Bin_OR = '0') then
         s_Energy_Bin_415 <= s_Energy_Bin_415 +'1';
		 Energy_Bin_Rdy_415 <= '1';
		else
		 s_Energy_Bin_415 <= s_Energy_Bin_415;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_415 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_415;  
 
  
  Energy_Bin_416 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_416   <=  (others =>'0');
		Energy_Bin_Rdy_416 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E416_C1_L and PEAK_C1 <= s_E416_C1_H and Bin_OR = '0') then
         s_Energy_Bin_416 <= s_Energy_Bin_416 +'1';
		 Energy_Bin_Rdy_416 <= '1';
		else
		 s_Energy_Bin_416 <= s_Energy_Bin_416;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_416 <= '0';
      end if;
    end if;
  end process  Energy_Bin_416;   
  
 Energy_Bin_417 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_417   <=  (others =>'0');
		Energy_Bin_Rdy_417 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E417_C1_L and PEAK_C1 <= s_E417_C1_H and Bin_OR = '0') then
         s_Energy_Bin_417 <= s_Energy_Bin_417 +'1';
		 Energy_Bin_Rdy_417 <= '1';
		else
		 s_Energy_Bin_417 <= s_Energy_Bin_417;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_417 <= '0';
      end if;
    end if;
  end process  Energy_Bin_417;   
  
  Energy_Bin_418 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_418   <=  (others =>'0');
		Energy_Bin_Rdy_418 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E418_C1_L and PEAK_C1 <= s_E418_C1_H and Bin_OR = '0') then
         s_Energy_Bin_418 <= s_Energy_Bin_418 +'1';
		 Energy_Bin_Rdy_418 <= '1';
		else
		 s_Energy_Bin_418 <= s_Energy_Bin_418;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_418 <= '0';
      end if;
    end if;
  end process  Energy_Bin_418;   
  
  Energy_Bin_419 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_419   <=  (others =>'0');
		Energy_Bin_Rdy_419 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E419_C1_L and PEAK_C1 <= s_E419_C1_H and Bin_OR = '0') then
         s_Energy_Bin_419 <= s_Energy_Bin_419 +'1';
		 Energy_Bin_Rdy_419 <= '1';
		else
		 s_Energy_Bin_419 <= s_Energy_Bin_419;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_419 <= '0';
      end if;
    end if;
  end process  Energy_Bin_419;       
  
     Energy_Bin_420 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_420   <=  (others =>'0');
		Energy_Bin_Rdy_420 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E420_C1_L and PEAK_C1 <= s_E420_C1_H and Bin_OR = '0') then
         s_Energy_Bin_420 <= s_Energy_Bin_420 +'1';
		 Energy_Bin_Rdy_420 <= '1';
		else
		 s_Energy_Bin_420 <= s_Energy_Bin_420;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_420 <= '0';
      end if;
    end if;
  end process  Energy_Bin_420;    
  
  Energy_Bin_421 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_421   <=  (others =>'0');
		Energy_Bin_Rdy_421 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E421_C1_L and PEAK_C1 <= s_E421_C1_H and Bin_OR = '0') then
         s_Energy_Bin_421 <= s_Energy_Bin_421 +'1';
		 Energy_Bin_Rdy_421 <= '1';
		else
		 s_Energy_Bin_421 <= s_Energy_Bin_421;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_421 <= '0';
      end if;
    end if;
  end process  Energy_Bin_421;   
  
  Energy_Bin_422 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_422   <=  (others =>'0');
	    Energy_Bin_Rdy_422 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E422_C1_L and PEAK_C1 <= s_E422_C1_H and Bin_OR = '0') then
         s_Energy_Bin_422 <= s_Energy_Bin_422 +'1';
		 Energy_Bin_Rdy_422 <= '1';
		else
		 s_Energy_Bin_422 <= s_Energy_Bin_422;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_422 <= '0';
      end if;
    end if;
  end process  Energy_Bin_422;   
  
  Energy_Bin_423 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_423   <=  (others =>'0');
	    Energy_Bin_Rdy_423 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E423_C1_L and PEAK_C1 <= s_E423_C1_H and Bin_OR = '0') then
         s_Energy_Bin_423 <= s_Energy_Bin_423 +'1';
		 Energy_Bin_Rdy_423 <= '1';
		else
		 s_Energy_Bin_423 <= s_Energy_Bin_423;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_423 <= '0';
      end if;
    end if;
  end process  Energy_Bin_423;   
  
  Energy_Bin_424 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_424   <=  (others =>'0');
		Energy_Bin_Rdy_424 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E424_C1_L and PEAK_C1 <= s_E424_C1_H and Bin_OR = '0') then
         s_Energy_Bin_424 <= s_Energy_Bin_424 +'1';
		 Energy_Bin_Rdy_424 <= '1';
		else
		 s_Energy_Bin_424 <= s_Energy_Bin_424;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_424 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_424;   
 
 
  Energy_Bin_425 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_425   <=  (others =>'0');
		Energy_Bin_Rdy_425 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E425_C1_L and PEAK_C1 <= s_E425_C1_H and Bin_OR = '0') then
         s_Energy_Bin_425 <= s_Energy_Bin_425 +'1';
		 Energy_Bin_Rdy_425 <= '1';
		else
		 s_Energy_Bin_425 <= s_Energy_Bin_425;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_425 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_425;  
 
  
  Energy_Bin_426 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_426   <=  (others =>'0');
		Energy_Bin_Rdy_426 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E426_C1_L and PEAK_C1 <= s_E426_C1_H and Bin_OR = '0') then
         s_Energy_Bin_426 <= s_Energy_Bin_426 +'1';
		 Energy_Bin_Rdy_426 <= '1';
		else
		 s_Energy_Bin_426 <= s_Energy_Bin_426;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_426 <= '0';
      end if;
    end if;
  end process  Energy_Bin_426;   
  
 Energy_Bin_427 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_427   <=  (others =>'0');
		Energy_Bin_Rdy_427 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E427_C1_L and PEAK_C1 <= s_E427_C1_H and Bin_OR = '0') then
         s_Energy_Bin_427 <= s_Energy_Bin_427 +'1';
		 Energy_Bin_Rdy_427 <= '1';
		else
		 s_Energy_Bin_427 <= s_Energy_Bin_427;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_427 <= '0';
      end if;
    end if;
  end process  Energy_Bin_427;   
  
  Energy_Bin_428 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_428   <=  (others =>'0');
		Energy_Bin_Rdy_428 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E428_C1_L and PEAK_C1 <= s_E428_C1_H and Bin_OR = '0') then
         s_Energy_Bin_428 <= s_Energy_Bin_428 +'1';
		 Energy_Bin_Rdy_428 <= '1';
		else
		 s_Energy_Bin_428 <= s_Energy_Bin_428;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_428 <= '0';
      end if;
    end if;
  end process  Energy_Bin_428;   
  
  Energy_Bin_429 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_429   <=  (others =>'0');
		Energy_Bin_Rdy_429 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E429_C1_L and PEAK_C1 <= s_E429_C1_H and Bin_OR = '0') then
         s_Energy_Bin_429 <= s_Energy_Bin_429 +'1';
		 Energy_Bin_Rdy_429 <= '1';
		else
		 s_Energy_Bin_429 <= s_Energy_Bin_429;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_429 <= '0';
      end if;
    end if;
  end process  Energy_Bin_429;        
  
     Energy_Bin_430 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_430   <=  (others =>'0');
		Energy_Bin_Rdy_430 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E430_C1_L and PEAK_C1 <= s_E430_C1_H and Bin_OR = '0') then
         s_Energy_Bin_430 <= s_Energy_Bin_430 +'1';
		 Energy_Bin_Rdy_430 <= '1';
		else
		 s_Energy_Bin_430 <= s_Energy_Bin_430;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_430 <= '0';
      end if;
    end if;
  end process  Energy_Bin_430;    
  
  Energy_Bin_431 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_431   <=  (others =>'0');
		Energy_Bin_Rdy_431 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E431_C1_L and PEAK_C1 <= s_E431_C1_H and Bin_OR = '0') then
         s_Energy_Bin_431 <= s_Energy_Bin_431 +'1';
		 Energy_Bin_Rdy_431 <= '1';
		else
		 s_Energy_Bin_431 <= s_Energy_Bin_431;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_431 <= '0';
      end if;
    end if;
  end process  Energy_Bin_431;   
  
  Energy_Bin_432 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_432   <=  (others =>'0');
	    Energy_Bin_Rdy_432 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E432_C1_L and PEAK_C1 <= s_E432_C1_H and Bin_OR = '0') then
         s_Energy_Bin_432 <= s_Energy_Bin_432 +'1';
		 Energy_Bin_Rdy_432 <= '1';
		else
		 s_Energy_Bin_432 <= s_Energy_Bin_432;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_432 <= '0';
      end if;
    end if;
  end process  Energy_Bin_432;   
  
  Energy_Bin_433 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_433   <=  (others =>'0');
	    Energy_Bin_Rdy_433 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E433_C1_L and PEAK_C1 <= s_E433_C1_H and Bin_OR = '0') then
         s_Energy_Bin_433 <= s_Energy_Bin_433 +'1';
		 Energy_Bin_Rdy_433 <= '1';
		else
		 s_Energy_Bin_433 <= s_Energy_Bin_433;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_433 <= '0';
      end if;
    end if;
  end process  Energy_Bin_433;   
  
  Energy_Bin_434 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_434   <=  (others =>'0');
		Energy_Bin_Rdy_434 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E434_C1_L and PEAK_C1 <= s_E434_C1_H and Bin_OR = '0') then
         s_Energy_Bin_434 <= s_Energy_Bin_434 +'1';
		 Energy_Bin_Rdy_434 <= '1';
		else
		 s_Energy_Bin_434 <= s_Energy_Bin_434;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_434 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_434;   
 
 
  Energy_Bin_435 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_435   <=  (others =>'0');
		Energy_Bin_Rdy_435 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E435_C1_L and PEAK_C1 <= s_E435_C1_H and Bin_OR = '0') then
         s_Energy_Bin_435 <= s_Energy_Bin_435 +'1';
		 Energy_Bin_Rdy_435 <= '1';
		else
		 s_Energy_Bin_435 <= s_Energy_Bin_435;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_435 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_435;  
 
  
  Energy_Bin_436 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_436   <=  (others =>'0');
		Energy_Bin_Rdy_436 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E436_C1_L and PEAK_C1 <= s_E436_C1_H and Bin_OR = '0') then
         s_Energy_Bin_436 <= s_Energy_Bin_436 +'1';
		 Energy_Bin_Rdy_436 <= '1';
		else
		 s_Energy_Bin_436 <= s_Energy_Bin_436;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_436 <= '0';
      end if;
    end if;
  end process  Energy_Bin_436;   
  
 Energy_Bin_437 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_437   <=  (others =>'0');
		Energy_Bin_Rdy_437 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E437_C1_L and PEAK_C1 <= s_E437_C1_H and Bin_OR = '0') then
         s_Energy_Bin_437 <= s_Energy_Bin_437 +'1';
		 Energy_Bin_Rdy_437 <= '1';
		else
		 s_Energy_Bin_437 <= s_Energy_Bin_437;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_437 <= '0';
      end if;
    end if;
  end process  Energy_Bin_437;   
  
  Energy_Bin_438 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_438   <=  (others =>'0');
		Energy_Bin_Rdy_438 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E438_C1_L and PEAK_C1 <= s_E438_C1_H and Bin_OR = '0') then
         s_Energy_Bin_438 <= s_Energy_Bin_438 +'1';
		 Energy_Bin_Rdy_438 <= '1';
		else
		 s_Energy_Bin_438 <= s_Energy_Bin_438;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_438 <= '0';
      end if;
    end if;
  end process  Energy_Bin_438;   
  
  Energy_Bin_439 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_439   <=  (others =>'0');
		Energy_Bin_Rdy_439 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E439_C1_L and PEAK_C1 <= s_E439_C1_H and Bin_OR = '0') then
         s_Energy_Bin_439 <= s_Energy_Bin_439 +'1';
		 Energy_Bin_Rdy_439 <= '1';
		else
		 s_Energy_Bin_439 <= s_Energy_Bin_439;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_439 <= '0';
      end if;
    end if;
  end process  Energy_Bin_439;         
  
     Energy_Bin_440 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_440   <=  (others =>'0');
		Energy_Bin_Rdy_440 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E440_C1_L and PEAK_C1 <= s_E440_C1_H and Bin_OR = '0') then
         s_Energy_Bin_440 <= s_Energy_Bin_440 +'1';
		 Energy_Bin_Rdy_440 <= '1';
		else
		 s_Energy_Bin_440 <= s_Energy_Bin_440;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_440 <= '0';
      end if;
    end if;
  end process  Energy_Bin_440;    
  
  Energy_Bin_441 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_441   <=  (others =>'0');
		Energy_Bin_Rdy_441 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E441_C1_L and PEAK_C1 <= s_E441_C1_H and Bin_OR = '0') then
         s_Energy_Bin_441 <= s_Energy_Bin_441 +'1';
		 Energy_Bin_Rdy_441 <= '1';
		else
		 s_Energy_Bin_441 <= s_Energy_Bin_441;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_441 <= '0';
      end if;
    end if;
  end process  Energy_Bin_441;   
  
  Energy_Bin_442 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_442   <=  (others =>'0');
	    Energy_Bin_Rdy_442 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E442_C1_L and PEAK_C1 <= s_E442_C1_H and Bin_OR = '0') then
         s_Energy_Bin_442 <= s_Energy_Bin_442 +'1';
		 Energy_Bin_Rdy_442 <= '1';
		else
		 s_Energy_Bin_442 <= s_Energy_Bin_442;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_442 <= '0';
      end if;
    end if;
  end process  Energy_Bin_442;   
  
  Energy_Bin_443 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_443   <=  (others =>'0');
	    Energy_Bin_Rdy_443 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E443_C1_L and PEAK_C1 <= s_E443_C1_H and Bin_OR = '0') then
         s_Energy_Bin_443 <= s_Energy_Bin_443 +'1';
		 Energy_Bin_Rdy_443 <= '1';
		else
		 s_Energy_Bin_443 <= s_Energy_Bin_443;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_443 <= '0';
      end if;
    end if;
  end process  Energy_Bin_443;   
  
  Energy_Bin_444 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_444   <=  (others =>'0');
		Energy_Bin_Rdy_444 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E444_C1_L and PEAK_C1 <= s_E444_C1_H and Bin_OR = '0') then
         s_Energy_Bin_444 <= s_Energy_Bin_444 +'1';
		 Energy_Bin_Rdy_444 <= '1';
		else
		 s_Energy_Bin_444 <= s_Energy_Bin_444;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_444 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_444;   
 
 
  Energy_Bin_445 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_445   <=  (others =>'0');
		Energy_Bin_Rdy_445 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E445_C1_L and PEAK_C1 <= s_E445_C1_H and Bin_OR = '0') then
         s_Energy_Bin_445 <= s_Energy_Bin_445 +'1';
		 Energy_Bin_Rdy_445 <= '1';
		else
		 s_Energy_Bin_445 <= s_Energy_Bin_445;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_445 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_445;  
 
  
  Energy_Bin_446 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_446   <=  (others =>'0');
		Energy_Bin_Rdy_446 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E446_C1_L and PEAK_C1 <= s_E446_C1_H and Bin_OR = '0') then
         s_Energy_Bin_446 <= s_Energy_Bin_446 +'1';
		 Energy_Bin_Rdy_446 <= '1';
		else
		 s_Energy_Bin_446 <= s_Energy_Bin_446;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_446 <= '0';
      end if;
    end if;
  end process  Energy_Bin_446;   
  
 Energy_Bin_447 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_447   <=  (others =>'0');
		Energy_Bin_Rdy_447 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E447_C1_L and PEAK_C1 <= s_E447_C1_H and Bin_OR = '0') then
         s_Energy_Bin_447 <= s_Energy_Bin_447 +'1';
		 Energy_Bin_Rdy_447 <= '1';
		else
		 s_Energy_Bin_447 <= s_Energy_Bin_447;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_447 <= '0';
      end if;
    end if;
  end process  Energy_Bin_447;   
  
  Energy_Bin_448 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_448   <=  (others =>'0');
		Energy_Bin_Rdy_448 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E448_C1_L and PEAK_C1 <= s_E448_C1_H and Bin_OR = '0') then
         s_Energy_Bin_448 <= s_Energy_Bin_448 +'1';
		 Energy_Bin_Rdy_448 <= '1';
		else
		 s_Energy_Bin_448 <= s_Energy_Bin_448;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_448 <= '0';
      end if;
    end if;
  end process  Energy_Bin_448;   
  
  Energy_Bin_449 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_449   <=  (others =>'0');
		Energy_Bin_Rdy_449 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E449_C1_L and PEAK_C1 <= s_E449_C1_H and Bin_OR = '0') then
         s_Energy_Bin_449 <= s_Energy_Bin_449 +'1';
		 Energy_Bin_Rdy_449 <= '1';
		else
		 s_Energy_Bin_449 <= s_Energy_Bin_449;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_449 <= '0';
      end if;
    end if;
  end process  Energy_Bin_449;          
  
  
     Energy_Bin_450 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_450   <=  (others =>'0');
		Energy_Bin_Rdy_450 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E450_C1_L and PEAK_C1 <= s_E450_C1_H and Bin_OR = '0') then
         s_Energy_Bin_450 <= s_Energy_Bin_450 +'1';
		 Energy_Bin_Rdy_450 <= '1';
		else
		 s_Energy_Bin_450 <= s_Energy_Bin_450;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_450 <= '0';
      end if;
    end if;
  end process  Energy_Bin_450;    
  
  Energy_Bin_451 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_451   <=  (others =>'0');
		Energy_Bin_Rdy_451 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E451_C1_L and PEAK_C1 <= s_E451_C1_H and Bin_OR = '0') then
         s_Energy_Bin_451 <= s_Energy_Bin_451 +'1';
		 Energy_Bin_Rdy_451 <= '1';
		else
		 s_Energy_Bin_451 <= s_Energy_Bin_451;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_451 <= '0';
      end if;
    end if;
  end process  Energy_Bin_451;   
  
  Energy_Bin_452 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_452   <=  (others =>'0');
	    Energy_Bin_Rdy_452 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E452_C1_L and PEAK_C1 <= s_E452_C1_H and Bin_OR = '0') then
         s_Energy_Bin_452 <= s_Energy_Bin_452 +'1';
		 Energy_Bin_Rdy_452 <= '1';
		else
		 s_Energy_Bin_452 <= s_Energy_Bin_452;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_452 <= '0';
      end if;
    end if;
  end process  Energy_Bin_452;   
  
  Energy_Bin_453 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_453   <=  (others =>'0');
	    Energy_Bin_Rdy_453 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E453_C1_L and PEAK_C1 <= s_E453_C1_H and Bin_OR = '0') then
         s_Energy_Bin_453 <= s_Energy_Bin_453 +'1';
		 Energy_Bin_Rdy_453 <= '1';
		else
		 s_Energy_Bin_453 <= s_Energy_Bin_453;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_453 <= '0';
      end if;
    end if;
  end process  Energy_Bin_453;   
  
  Energy_Bin_454 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_454   <=  (others =>'0');
		Energy_Bin_Rdy_454 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E454_C1_L and PEAK_C1 <= s_E454_C1_H and Bin_OR = '0') then
         s_Energy_Bin_454 <= s_Energy_Bin_454 +'1';
		 Energy_Bin_Rdy_454 <= '1';
		else
		 s_Energy_Bin_454 <= s_Energy_Bin_454;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_454 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_454;   
 
 
  Energy_Bin_455 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_455   <=  (others =>'0');
		Energy_Bin_Rdy_455 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E455_C1_L and PEAK_C1 <= s_E455_C1_H and Bin_OR = '0') then
         s_Energy_Bin_455 <= s_Energy_Bin_455 +'1';
		 Energy_Bin_Rdy_455 <= '1';
		else
		 s_Energy_Bin_455 <= s_Energy_Bin_455;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_455 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_455;  
 
  
  Energy_Bin_456 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_456   <=  (others =>'0');
		Energy_Bin_Rdy_456 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E456_C1_L and PEAK_C1 <= s_E456_C1_H and Bin_OR = '0') then
         s_Energy_Bin_456 <= s_Energy_Bin_456 +'1';
		 Energy_Bin_Rdy_456 <= '1';
		else
		 s_Energy_Bin_456 <= s_Energy_Bin_456;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_456 <= '0';
      end if;
    end if;
  end process  Energy_Bin_456;   
  
 Energy_Bin_457 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_457   <=  (others =>'0');
		Energy_Bin_Rdy_457 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E457_C1_L and PEAK_C1 <= s_E457_C1_H and Bin_OR = '0') then
         s_Energy_Bin_457 <= s_Energy_Bin_457 +'1';
		 Energy_Bin_Rdy_457 <= '1';
		else
		 s_Energy_Bin_457 <= s_Energy_Bin_457;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_457 <= '0';
      end if;
    end if;
  end process  Energy_Bin_457;   
  
  Energy_Bin_458 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_458   <=  (others =>'0');
		Energy_Bin_Rdy_458 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E458_C1_L and PEAK_C1 <= s_E458_C1_H and Bin_OR = '0') then
         s_Energy_Bin_458 <= s_Energy_Bin_458 +'1';
		 Energy_Bin_Rdy_458 <= '1';
		else
		 s_Energy_Bin_458 <= s_Energy_Bin_458;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_458 <= '0';
      end if;
    end if;
  end process  Energy_Bin_458;   
  
  Energy_Bin_459 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_459   <=  (others =>'0');
		Energy_Bin_Rdy_459 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E459_C1_L and PEAK_C1 <= s_E459_C1_H and Bin_OR = '0') then
         s_Energy_Bin_459 <= s_Energy_Bin_459 +'1';
		 Energy_Bin_Rdy_459 <= '1';
		else
		 s_Energy_Bin_459 <= s_Energy_Bin_459;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_459 <= '0';
      end if;
    end if;
  end process  Energy_Bin_459;           
  
     Energy_Bin_460 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_460   <=  (others =>'0');
		Energy_Bin_Rdy_460 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E460_C1_L and PEAK_C1 <= s_E460_C1_H and Bin_OR = '0') then
         s_Energy_Bin_460 <= s_Energy_Bin_460 +'1';
		 Energy_Bin_Rdy_460 <= '1';
		else
		 s_Energy_Bin_460 <= s_Energy_Bin_460;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_460 <= '0';
      end if;
    end if;
  end process  Energy_Bin_460;    
  
  Energy_Bin_461 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_461   <=  (others =>'0');
		Energy_Bin_Rdy_461 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E461_C1_L and PEAK_C1 <= s_E461_C1_H and Bin_OR = '0') then
         s_Energy_Bin_461 <= s_Energy_Bin_461 +'1';
		 Energy_Bin_Rdy_461 <= '1';
		else
		 s_Energy_Bin_461 <= s_Energy_Bin_461;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_461 <= '0';
      end if;
    end if;
  end process  Energy_Bin_461;   
  
  Energy_Bin_462 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_462   <=  (others =>'0');
	    Energy_Bin_Rdy_462 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E462_C1_L and PEAK_C1 <= s_E462_C1_H and Bin_OR = '0') then
         s_Energy_Bin_462 <= s_Energy_Bin_462 +'1';
		 Energy_Bin_Rdy_462 <= '1';
		else
		 s_Energy_Bin_462 <= s_Energy_Bin_462;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_462 <= '0';
      end if;
    end if;
  end process  Energy_Bin_462;   
  
  Energy_Bin_463 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_463   <=  (others =>'0');
	    Energy_Bin_Rdy_463 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E463_C1_L and PEAK_C1 <= s_E463_C1_H and Bin_OR = '0') then
         s_Energy_Bin_463 <= s_Energy_Bin_463 +'1';
		 Energy_Bin_Rdy_463 <= '1';
		else
		 s_Energy_Bin_463 <= s_Energy_Bin_463;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_463 <= '0';
      end if;
    end if;
  end process  Energy_Bin_463;   
  
  Energy_Bin_464 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_464   <=  (others =>'0');
		Energy_Bin_Rdy_464 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E464_C1_L and PEAK_C1 <= s_E464_C1_H and Bin_OR = '0') then
         s_Energy_Bin_464 <= s_Energy_Bin_464 +'1';
		 Energy_Bin_Rdy_464 <= '1';
		else
		 s_Energy_Bin_464 <= s_Energy_Bin_464;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_464 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_464;   
 
 
  Energy_Bin_465 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_465   <=  (others =>'0');
		Energy_Bin_Rdy_465 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E465_C1_L and PEAK_C1 <= s_E465_C1_H and Bin_OR = '0') then
         s_Energy_Bin_465 <= s_Energy_Bin_465 +'1';
		 Energy_Bin_Rdy_465 <= '1';
		else
		 s_Energy_Bin_465 <= s_Energy_Bin_465;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_465 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_465;  
 
  
  Energy_Bin_466 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_466   <=  (others =>'0');
		Energy_Bin_Rdy_466 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E466_C1_L and PEAK_C1 <= s_E466_C1_H and Bin_OR = '0') then
         s_Energy_Bin_466 <= s_Energy_Bin_466 +'1';
		 Energy_Bin_Rdy_466 <= '1';
		else
		 s_Energy_Bin_466 <= s_Energy_Bin_466;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_466 <= '0';
      end if;
    end if;
  end process  Energy_Bin_466;   
  
 Energy_Bin_467 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_467   <=  (others =>'0');
		Energy_Bin_Rdy_467 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E467_C1_L and PEAK_C1 <= s_E467_C1_H and Bin_OR = '0') then
         s_Energy_Bin_467 <= s_Energy_Bin_467 +'1';
		 Energy_Bin_Rdy_467 <= '1';
		else
		 s_Energy_Bin_467 <= s_Energy_Bin_467;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_467 <= '0';
      end if;
    end if;
  end process  Energy_Bin_467;   
  
  Energy_Bin_468 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_468   <=  (others =>'0');
		Energy_Bin_Rdy_468 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E468_C1_L and PEAK_C1 <= s_E468_C1_H and Bin_OR = '0') then
         s_Energy_Bin_468 <= s_Energy_Bin_468 +'1';
		 Energy_Bin_Rdy_468 <= '1';
		else
		 s_Energy_Bin_468 <= s_Energy_Bin_468;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_468 <= '0';
      end if;
    end if;
  end process  Energy_Bin_468;   
  
  Energy_Bin_469 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_469   <=  (others =>'0');
		Energy_Bin_Rdy_469 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E469_C1_L and PEAK_C1 <= s_E469_C1_H and Bin_OR = '0') then
         s_Energy_Bin_469 <= s_Energy_Bin_469 +'1';
		 Energy_Bin_Rdy_469 <= '1';
		else
		 s_Energy_Bin_469 <= s_Energy_Bin_469;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_469 <= '0';
      end if;
    end if;
  end process  Energy_Bin_469;         
  
     Energy_Bin_470 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_470   <=  (others =>'0');
		Energy_Bin_Rdy_470 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E470_C1_L and PEAK_C1 <= s_E470_C1_H and Bin_OR = '0') then
         s_Energy_Bin_470 <= s_Energy_Bin_470 +'1';
		 Energy_Bin_Rdy_470 <= '1';
		else
		 s_Energy_Bin_470 <= s_Energy_Bin_470;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_470 <= '0';
      end if;
    end if;
  end process  Energy_Bin_470;    
  
  Energy_Bin_471 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_471   <=  (others =>'0');
		Energy_Bin_Rdy_471 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E471_C1_L and PEAK_C1 <= s_E471_C1_H and Bin_OR = '0') then
         s_Energy_Bin_471 <= s_Energy_Bin_471 +'1';
		 Energy_Bin_Rdy_471 <= '1';
		else
		 s_Energy_Bin_471 <= s_Energy_Bin_471;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_471 <= '0';
      end if;
    end if;
  end process  Energy_Bin_471;   
  
  Energy_Bin_472 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_472   <=  (others =>'0');
	    Energy_Bin_Rdy_472 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E472_C1_L and PEAK_C1 <= s_E472_C1_H and Bin_OR = '0') then
         s_Energy_Bin_472 <= s_Energy_Bin_472 +'1';
		 Energy_Bin_Rdy_472 <= '1';
		else
		 s_Energy_Bin_472 <= s_Energy_Bin_472;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_472 <= '0';
      end if;
    end if;
  end process  Energy_Bin_472;   
  
  Energy_Bin_473 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_473   <=  (others =>'0');
	    Energy_Bin_Rdy_473 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E473_C1_L and PEAK_C1 <= s_E473_C1_H and Bin_OR = '0') then
         s_Energy_Bin_473 <= s_Energy_Bin_473 +'1';
		 Energy_Bin_Rdy_473 <= '1';
		else
		 s_Energy_Bin_473 <= s_Energy_Bin_473;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_473 <= '0';
      end if;
    end if;
  end process  Energy_Bin_473;   
  
  Energy_Bin_474 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_474   <=  (others =>'0');
		Energy_Bin_Rdy_474 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E474_C1_L and PEAK_C1 <= s_E474_C1_H and Bin_OR = '0') then
         s_Energy_Bin_474 <= s_Energy_Bin_474 +'1';
		 Energy_Bin_Rdy_474 <= '1';
		else
		 s_Energy_Bin_474 <= s_Energy_Bin_474;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_474 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_474;   
 
 
  Energy_Bin_475 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_475   <=  (others =>'0');
		Energy_Bin_Rdy_475 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E475_C1_L and PEAK_C1 <= s_E475_C1_H and Bin_OR = '0') then
         s_Energy_Bin_475 <= s_Energy_Bin_475 +'1';
		 Energy_Bin_Rdy_475 <= '1';
		else
		 s_Energy_Bin_475 <= s_Energy_Bin_475;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_475 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_475;  
 
  
  Energy_Bin_476 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_476   <=  (others =>'0');
		Energy_Bin_Rdy_476 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E476_C1_L and PEAK_C1 <= s_E476_C1_H and Bin_OR = '0') then
         s_Energy_Bin_476 <= s_Energy_Bin_476 +'1';
		 Energy_Bin_Rdy_476 <= '1';
		else
		 s_Energy_Bin_476 <= s_Energy_Bin_476;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_476 <= '0';
      end if;
    end if;
  end process  Energy_Bin_476;   
  
 Energy_Bin_477 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_477   <=  (others =>'0');
		Energy_Bin_Rdy_477 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E477_C1_L and PEAK_C1 <= s_E477_C1_H and Bin_OR = '0') then
         s_Energy_Bin_477 <= s_Energy_Bin_477 +'1';
		 Energy_Bin_Rdy_477 <= '1';
		else
		 s_Energy_Bin_477 <= s_Energy_Bin_477;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_477 <= '0';
      end if;
    end if;
  end process  Energy_Bin_477;   
  
  Energy_Bin_478 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_478   <=  (others =>'0');
		Energy_Bin_Rdy_478 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E478_C1_L and PEAK_C1 <= s_E478_C1_H and Bin_OR = '0') then
         s_Energy_Bin_478 <= s_Energy_Bin_478 +'1';
		 Energy_Bin_Rdy_478 <= '1';
		else
		 s_Energy_Bin_478 <= s_Energy_Bin_478;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_478 <= '0';
      end if;
    end if;
  end process  Energy_Bin_478;   
  
  Energy_Bin_479 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_479   <=  (others =>'0');
		Energy_Bin_Rdy_479 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E479_C1_L and PEAK_C1 <= s_E479_C1_H and Bin_OR = '0') then
         s_Energy_Bin_479 <= s_Energy_Bin_479 +'1';
		 Energy_Bin_Rdy_479 <= '1';
		else
		 s_Energy_Bin_479 <= s_Energy_Bin_479;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_479 <= '0';
      end if;
    end if;
  end process  Energy_Bin_479;       
  
     Energy_Bin_480 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_480   <=  (others =>'0');
		Energy_Bin_Rdy_480 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E480_C1_L and PEAK_C1 <= s_E480_C1_H and Bin_OR = '0') then
         s_Energy_Bin_480 <= s_Energy_Bin_480 +'1';
		 Energy_Bin_Rdy_480 <= '1';
		else
		 s_Energy_Bin_480 <= s_Energy_Bin_480;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_480 <= '0';
      end if;
    end if;
  end process  Energy_Bin_480;    
  
  Energy_Bin_481 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_481   <=  (others =>'0');
		Energy_Bin_Rdy_481 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E481_C1_L and PEAK_C1 <= s_E481_C1_H and Bin_OR = '0') then
         s_Energy_Bin_481 <= s_Energy_Bin_481 +'1';
		 Energy_Bin_Rdy_481 <= '1';
		else
		 s_Energy_Bin_481 <= s_Energy_Bin_481;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_481 <= '0';
      end if;
    end if;
  end process  Energy_Bin_481;   
  
  Energy_Bin_482 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_482   <=  (others =>'0');
	    Energy_Bin_Rdy_482 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E482_C1_L and PEAK_C1 <= s_E482_C1_H and Bin_OR = '0') then
         s_Energy_Bin_482 <= s_Energy_Bin_482 +'1';
		 Energy_Bin_Rdy_482 <= '1';
		else
		 s_Energy_Bin_482 <= s_Energy_Bin_482;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_482 <= '0';
      end if;
    end if;
  end process  Energy_Bin_482;   
  
  Energy_Bin_483 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_483   <=  (others =>'0');
	    Energy_Bin_Rdy_483 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E483_C1_L and PEAK_C1 <= s_E483_C1_H and Bin_OR = '0') then
         s_Energy_Bin_483 <= s_Energy_Bin_483 +'1';
		 Energy_Bin_Rdy_483 <= '1';
		else
		 s_Energy_Bin_483 <= s_Energy_Bin_483;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_483 <= '0';
      end if;
    end if;
  end process  Energy_Bin_483;   
  
  Energy_Bin_484 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_484   <=  (others =>'0');
		Energy_Bin_Rdy_484 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E484_C1_L and PEAK_C1 <= s_E484_C1_H and Bin_OR = '0') then
         s_Energy_Bin_484 <= s_Energy_Bin_484 +'1';
		 Energy_Bin_Rdy_484 <= '1';
		else
		 s_Energy_Bin_484 <= s_Energy_Bin_484;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_484 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_484;   
 
 
  Energy_Bin_485 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_485   <=  (others =>'0');
		Energy_Bin_Rdy_485 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E485_C1_L and PEAK_C1 <= s_E485_C1_H and Bin_OR = '0') then
         s_Energy_Bin_485 <= s_Energy_Bin_485 +'1';
		 Energy_Bin_Rdy_485 <= '1';
		else
		 s_Energy_Bin_485 <= s_Energy_Bin_485;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_485 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_485;  
 
  
  Energy_Bin_486 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_486   <=  (others =>'0');
		Energy_Bin_Rdy_486 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E486_C1_L and PEAK_C1 <= s_E486_C1_H and Bin_OR = '0') then
         s_Energy_Bin_486 <= s_Energy_Bin_486 +'1';
		 Energy_Bin_Rdy_486 <= '1';
		else
		 s_Energy_Bin_486 <= s_Energy_Bin_486;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_486 <= '0';
      end if;
    end if;
  end process  Energy_Bin_486;   
  
 Energy_Bin_487 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_487   <=  (others =>'0');
		Energy_Bin_Rdy_487 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E487_C1_L and PEAK_C1 <= s_E487_C1_H and Bin_OR = '0') then
         s_Energy_Bin_487 <= s_Energy_Bin_487 +'1';
		 Energy_Bin_Rdy_487 <= '1';
		else
		 s_Energy_Bin_487 <= s_Energy_Bin_487;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_487 <= '0';
      end if;
    end if;
  end process  Energy_Bin_487;   
  
  Energy_Bin_488 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_488   <=  (others =>'0');
		Energy_Bin_Rdy_488 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E488_C1_L and PEAK_C1 <= s_E488_C1_H and Bin_OR = '0') then
         s_Energy_Bin_488 <= s_Energy_Bin_488 +'1';
		 Energy_Bin_Rdy_488 <= '1';
		else
		 s_Energy_Bin_488 <= s_Energy_Bin_488;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_488 <= '0';
      end if;
    end if;
  end process  Energy_Bin_488;   
  
  Energy_Bin_489 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_489   <=  (others =>'0');
		Energy_Bin_Rdy_489 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E489_C1_L and PEAK_C1 <= s_E489_C1_H and Bin_OR = '0') then
         s_Energy_Bin_489 <= s_Energy_Bin_489 +'1';
		 Energy_Bin_Rdy_489 <= '1';
		else
		 s_Energy_Bin_489 <= s_Energy_Bin_489;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_489 <= '0';
      end if;
    end if;
  end process  Energy_Bin_489;      
  
     Energy_Bin_490 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_490   <=  (others =>'0');
		Energy_Bin_Rdy_490 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E490_C1_L and PEAK_C1 <= s_E490_C1_H and Bin_OR = '0') then
         s_Energy_Bin_490 <= s_Energy_Bin_490 +'1';
		 Energy_Bin_Rdy_490 <= '1';
		else
		 s_Energy_Bin_490 <= s_Energy_Bin_490;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_490 <= '0';
      end if;
    end if;
  end process  Energy_Bin_490;    
  
  Energy_Bin_491 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_491   <=  (others =>'0');
		Energy_Bin_Rdy_491 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E491_C1_L and PEAK_C1 <= s_E491_C1_H and Bin_OR = '0') then
         s_Energy_Bin_491 <= s_Energy_Bin_491 +'1';
		 Energy_Bin_Rdy_491 <= '1';
		else
		 s_Energy_Bin_491 <= s_Energy_Bin_491;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_491 <= '0';
      end if;
    end if;
  end process  Energy_Bin_491;   
  
  Energy_Bin_492 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_492   <=  (others =>'0');
	    Energy_Bin_Rdy_492 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E492_C1_L and PEAK_C1 <= s_E492_C1_H and Bin_OR = '0') then
         s_Energy_Bin_492 <= s_Energy_Bin_492 +'1';
		 Energy_Bin_Rdy_492 <= '1';
		else
		 s_Energy_Bin_492 <= s_Energy_Bin_492;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_492 <= '0';
      end if;
    end if;
  end process  Energy_Bin_492;   
  
  Energy_Bin_493 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_493   <=  (others =>'0');
	    Energy_Bin_Rdy_493 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E493_C1_L and PEAK_C1 <= s_E493_C1_H and Bin_OR = '0') then
         s_Energy_Bin_493 <= s_Energy_Bin_493 +'1';
		 Energy_Bin_Rdy_493 <= '1';
		else
		 s_Energy_Bin_493 <= s_Energy_Bin_493;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_493 <= '0';
      end if;
    end if;
  end process  Energy_Bin_493;   
  
  Energy_Bin_494 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_494   <=  (others =>'0');
		Energy_Bin_Rdy_494 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E494_C1_L and PEAK_C1 <= s_E494_C1_H and Bin_OR = '0') then
         s_Energy_Bin_494 <= s_Energy_Bin_494 +'1';
		 Energy_Bin_Rdy_494 <= '1';
		else
		 s_Energy_Bin_494 <= s_Energy_Bin_494;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_494 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_494;   
 
 
  Energy_Bin_495 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_495   <=  (others =>'0');
		Energy_Bin_Rdy_495 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E495_C1_L and PEAK_C1 <= s_E495_C1_H and Bin_OR = '0') then
         s_Energy_Bin_495 <= s_Energy_Bin_495 +'1';
		 Energy_Bin_Rdy_495 <= '1';
		else
		 s_Energy_Bin_495 <= s_Energy_Bin_495;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_495 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_495;  
 
  
  Energy_Bin_496 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_496   <=  (others =>'0');
		Energy_Bin_Rdy_496 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E496_C1_L and PEAK_C1 <= s_E496_C1_H and Bin_OR = '0') then
         s_Energy_Bin_496 <= s_Energy_Bin_496 +'1';
		 Energy_Bin_Rdy_496 <= '1';
		else
		 s_Energy_Bin_496 <= s_Energy_Bin_496;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_496 <= '0';
      end if;
    end if;
  end process  Energy_Bin_496;   
  
 Energy_Bin_497 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_497   <=  (others =>'0');
		Energy_Bin_Rdy_497 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E497_C1_L and PEAK_C1 <= s_E497_C1_H and Bin_OR = '0') then
         s_Energy_Bin_497 <= s_Energy_Bin_497 +'1';
		 Energy_Bin_Rdy_497 <= '1';
		else
		 s_Energy_Bin_497 <= s_Energy_Bin_497;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_497 <= '0';
      end if;
    end if;
  end process  Energy_Bin_497;   
  
  Energy_Bin_498 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_498   <=  (others =>'0');
		Energy_Bin_Rdy_498 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E498_C1_L and PEAK_C1 <= s_E498_C1_H and Bin_OR = '0') then
         s_Energy_Bin_498 <= s_Energy_Bin_498 +'1';
		 Energy_Bin_Rdy_498 <= '1';
		else
		 s_Energy_Bin_498 <= s_Energy_Bin_498;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_498 <= '0';
      end if;
    end if;
  end process  Energy_Bin_498;   
  
  Energy_Bin_499 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_499   <=  (others =>'0');
		Energy_Bin_Rdy_499 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E499_C1_L and PEAK_C1 <= s_E499_C1_H and Bin_OR = '0') then
         s_Energy_Bin_499 <= s_Energy_Bin_499 +'1';
		 Energy_Bin_Rdy_499 <= '1';
		else
		 s_Energy_Bin_499 <= s_Energy_Bin_499;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_499 <= '0';
      end if;
    end if;
  end process  Energy_Bin_499;      

    Energy_Bin_500 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_500   <=  (others =>'0');
		Energy_Bin_Rdy_500 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E500_C1_L and PEAK_C1 <= s_E500_C1_H and Bin_OR = '0') then
         s_Energy_Bin_500 <= s_Energy_Bin_500 +'1';
		 Energy_Bin_Rdy_500 <= '1';
		else
		 s_Energy_Bin_500 <= s_Energy_Bin_500;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_500 <= '0';
      end if;
    end if;
  end process  Energy_Bin_500;    
  
  Energy_Bin_501 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_501   <=  (others =>'0');
		Energy_Bin_Rdy_501 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E501_C1_L and PEAK_C1 <= s_E501_C1_H and Bin_OR = '0') then
         s_Energy_Bin_501 <= s_Energy_Bin_501 +'1';
		 Energy_Bin_Rdy_501 <= '1';
		else
		 s_Energy_Bin_501 <= s_Energy_Bin_501;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_501 <= '0';
      end if;
    end if;
  end process  Energy_Bin_501;   
  
  Energy_Bin_502 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_502   <=  (others =>'0');
	    Energy_Bin_Rdy_502 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E502_C1_L and PEAK_C1 <= s_E502_C1_H and Bin_OR = '0') then
         s_Energy_Bin_502 <= s_Energy_Bin_502 +'1';
		 Energy_Bin_Rdy_502 <= '1';
		else
		 s_Energy_Bin_502 <= s_Energy_Bin_502;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_502 <= '0';
      end if;
    end if;
  end process  Energy_Bin_502;   
  
  Energy_Bin_503 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_503   <=  (others =>'0');
	    Energy_Bin_Rdy_503 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E503_C1_L and PEAK_C1 <= s_E503_C1_H and Bin_OR = '0') then
         s_Energy_Bin_503 <= s_Energy_Bin_503 +'1';
		 Energy_Bin_Rdy_503 <= '1';
		else
		 s_Energy_Bin_503 <= s_Energy_Bin_503;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_503 <= '0';
      end if;
    end if;
  end process  Energy_Bin_503;   
  
  Energy_Bin_504 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_504   <=  (others =>'0');
		Energy_Bin_Rdy_504 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E504_C1_L and PEAK_C1 <= s_E504_C1_H and Bin_OR = '0') then
         s_Energy_Bin_504 <= s_Energy_Bin_504 +'1';
		 Energy_Bin_Rdy_504 <= '1';
		else
		 s_Energy_Bin_504 <= s_Energy_Bin_504;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_504 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_504;   
 
 
  Energy_Bin_505 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_505   <=  (others =>'0');
		Energy_Bin_Rdy_505 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E505_C1_L and PEAK_C1 <= s_E505_C1_H and Bin_OR = '0') then
         s_Energy_Bin_505 <= s_Energy_Bin_505 +'1';
		 Energy_Bin_Rdy_505 <= '1';
		else
		 s_Energy_Bin_505 <= s_Energy_Bin_505;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_505 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_505;  
 
  
  Energy_Bin_506 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_506   <=  (others =>'0');
		Energy_Bin_Rdy_506 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E506_C1_L and PEAK_C1 <= s_E506_C1_H and Bin_OR = '0') then
         s_Energy_Bin_506 <= s_Energy_Bin_506 +'1';
		 Energy_Bin_Rdy_506 <= '1';
		else
		 s_Energy_Bin_506 <= s_Energy_Bin_506;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_506 <= '0';
      end if;
    end if;
  end process  Energy_Bin_506;   
  
 Energy_Bin_507 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_507   <=  (others =>'0');
		Energy_Bin_Rdy_507 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E507_C1_L and PEAK_C1 <= s_E507_C1_H and Bin_OR = '0') then
         s_Energy_Bin_507 <= s_Energy_Bin_507 +'1';
		 Energy_Bin_Rdy_507 <= '1';
		else
		 s_Energy_Bin_507 <= s_Energy_Bin_507;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_507 <= '0';
      end if;
    end if;
  end process  Energy_Bin_507;   
  
  Energy_Bin_508 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_508   <=  (others =>'0');
		Energy_Bin_Rdy_508 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E508_C1_L and PEAK_C1 <= s_E508_C1_H and Bin_OR = '0') then
         s_Energy_Bin_508 <= s_Energy_Bin_508 +'1';
		 Energy_Bin_Rdy_508 <= '1';
		else
		 s_Energy_Bin_508 <= s_Energy_Bin_508;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_508 <= '0';
      end if;
    end if;
  end process  Energy_Bin_508;   
  
  Energy_Bin_509 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_509   <=  (others =>'0');
		Energy_Bin_Rdy_509 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E509_C1_L and PEAK_C1 <= s_E509_C1_H and Bin_OR = '0') then
         s_Energy_Bin_509 <= s_Energy_Bin_509 +'1';
		 Energy_Bin_Rdy_509 <= '1';
		else
		 s_Energy_Bin_509 <= s_Energy_Bin_509;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_509 <= '0';
      end if;
    end if;
  end process  Energy_Bin_509;      
  
     Energy_Bin_510 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_510   <=  (others =>'0');
		Energy_Bin_Rdy_510 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E510_C1_L and PEAK_C1 <= s_E510_C1_H and Bin_OR = '0') then
         s_Energy_Bin_510 <= s_Energy_Bin_510 +'1';
		 Energy_Bin_Rdy_510 <= '1';
		else
		 s_Energy_Bin_510 <= s_Energy_Bin_510;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_510 <= '0';
      end if;
    end if;
  end process  Energy_Bin_510;    
  
  Energy_Bin_511 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_511   <=  (others =>'0');
		Energy_Bin_Rdy_511 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E511_C1_L and PEAK_C1 <= s_E511_C1_H and Bin_OR = '0') then
         s_Energy_Bin_511 <= s_Energy_Bin_511 +'1';
		 Energy_Bin_Rdy_511 <= '1';
		else
		 s_Energy_Bin_511 <= s_Energy_Bin_511;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_511 <= '0';
      end if;
    end if;
  end process  Energy_Bin_511;   
  
  Energy_Bin_512 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_512   <=  (others =>'0');
	    Energy_Bin_Rdy_512 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E512_C1_L and PEAK_C1 <= s_E512_C1_H and Bin_OR = '0') then
         s_Energy_Bin_512 <= s_Energy_Bin_512 +'1';
		 Energy_Bin_Rdy_512 <= '1';
		else
		 s_Energy_Bin_512 <= s_Energy_Bin_512;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_512 <= '0';
      end if;
    end if;
  end process  Energy_Bin_512;   
  
  Energy_Bin_513 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_513   <=  (others =>'0');
	    Energy_Bin_Rdy_513 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E513_C1_L and PEAK_C1 <= s_E513_C1_H and Bin_OR = '0') then
         s_Energy_Bin_513 <= s_Energy_Bin_513 +'1';
		 Energy_Bin_Rdy_513 <= '1';
		else
		 s_Energy_Bin_513 <= s_Energy_Bin_513;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_513 <= '0';
      end if;
    end if;
  end process  Energy_Bin_513;   
  
  Energy_Bin_514 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_514   <=  (others =>'0');
		Energy_Bin_Rdy_514 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E514_C1_L and PEAK_C1 <= s_E514_C1_H and Bin_OR = '0') then
         s_Energy_Bin_514 <= s_Energy_Bin_514 +'1';
		 Energy_Bin_Rdy_514 <= '1';
		else
		 s_Energy_Bin_514 <= s_Energy_Bin_514;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_514 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_514;   
 
 
  Energy_Bin_515 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_515   <=  (others =>'0');
		Energy_Bin_Rdy_515 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E515_C1_L and PEAK_C1 <= s_E515_C1_H and Bin_OR = '0') then
         s_Energy_Bin_515 <= s_Energy_Bin_515 +'1';
		 Energy_Bin_Rdy_515 <= '1';
		else
		 s_Energy_Bin_515 <= s_Energy_Bin_515;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_515 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_515;  
 
  
  Energy_Bin_516 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_516   <=  (others =>'0');
		Energy_Bin_Rdy_516 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E516_C1_L and PEAK_C1 <= s_E516_C1_H and Bin_OR = '0') then
         s_Energy_Bin_516 <= s_Energy_Bin_516 +'1';
		 Energy_Bin_Rdy_516 <= '1';
		else
		 s_Energy_Bin_516 <= s_Energy_Bin_516;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_516 <= '0';
      end if;
    end if;
  end process  Energy_Bin_516;   
  
 Energy_Bin_517 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_517   <=  (others =>'0');
		Energy_Bin_Rdy_517 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E517_C1_L and PEAK_C1 <= s_E517_C1_H and Bin_OR = '0') then
         s_Energy_Bin_517 <= s_Energy_Bin_517 +'1';
		 Energy_Bin_Rdy_517 <= '1';
		else
		 s_Energy_Bin_517 <= s_Energy_Bin_517;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_517 <= '0';
      end if;
    end if;
  end process  Energy_Bin_517;   
  
  Energy_Bin_518 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_518   <=  (others =>'0');
		Energy_Bin_Rdy_518 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E518_C1_L and PEAK_C1 <= s_E518_C1_H and Bin_OR = '0') then
         s_Energy_Bin_518 <= s_Energy_Bin_518 +'1';
		 Energy_Bin_Rdy_518 <= '1';
		else
		 s_Energy_Bin_518 <= s_Energy_Bin_518;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_518 <= '0';
      end if;
    end if;
  end process  Energy_Bin_518;   
  
  Energy_Bin_519 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_519   <=  (others =>'0');
		Energy_Bin_Rdy_519 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E519_C1_L and PEAK_C1 <= s_E519_C1_H and Bin_OR = '0') then
         s_Energy_Bin_519 <= s_Energy_Bin_519 +'1';
		 Energy_Bin_Rdy_519 <= '1';
		else
		 s_Energy_Bin_519 <= s_Energy_Bin_519;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_519 <= '0';
      end if;
    end if;
  end process  Energy_Bin_519;       
  
     Energy_Bin_520 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_520   <=  (others =>'0');
		Energy_Bin_Rdy_520 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E520_C1_L and PEAK_C1 <= s_E520_C1_H and Bin_OR = '0') then
         s_Energy_Bin_520 <= s_Energy_Bin_520 +'1';
		 Energy_Bin_Rdy_520 <= '1';
		else
		 s_Energy_Bin_520 <= s_Energy_Bin_520;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_520 <= '0';
      end if;
    end if;
  end process  Energy_Bin_520;    
  
  Energy_Bin_521 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_521   <=  (others =>'0');
		Energy_Bin_Rdy_521 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E521_C1_L and PEAK_C1 <= s_E521_C1_H and Bin_OR = '0') then
         s_Energy_Bin_521 <= s_Energy_Bin_521 +'1';
		 Energy_Bin_Rdy_521 <= '1';
		else
		 s_Energy_Bin_521 <= s_Energy_Bin_521;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_521 <= '0';
      end if;
    end if;
  end process  Energy_Bin_521;   
  
  Energy_Bin_522 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_522   <=  (others =>'0');
	    Energy_Bin_Rdy_522 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E522_C1_L and PEAK_C1 <= s_E522_C1_H and Bin_OR = '0') then
         s_Energy_Bin_522 <= s_Energy_Bin_522 +'1';
		 Energy_Bin_Rdy_522 <= '1';
		else
		 s_Energy_Bin_522 <= s_Energy_Bin_522;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_522 <= '0';
      end if;
    end if;
  end process  Energy_Bin_522;   
  
  Energy_Bin_523 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_523   <=  (others =>'0');
	    Energy_Bin_Rdy_523 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E523_C1_L and PEAK_C1 <= s_E523_C1_H and Bin_OR = '0') then
         s_Energy_Bin_523 <= s_Energy_Bin_523 +'1';
		 Energy_Bin_Rdy_523 <= '1';
		else
		 s_Energy_Bin_523 <= s_Energy_Bin_523;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_523 <= '0';
      end if;
    end if;
  end process  Energy_Bin_523;   
  
  Energy_Bin_524 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_524   <=  (others =>'0');
		Energy_Bin_Rdy_524 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E524_C1_L and PEAK_C1 <= s_E524_C1_H and Bin_OR = '0') then
         s_Energy_Bin_524 <= s_Energy_Bin_524 +'1';
		 Energy_Bin_Rdy_524 <= '1';
		else
		 s_Energy_Bin_524 <= s_Energy_Bin_524;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_524 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_524;   
 
 
  Energy_Bin_525 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_525   <=  (others =>'0');
		Energy_Bin_Rdy_525 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E525_C1_L and PEAK_C1 <= s_E525_C1_H and Bin_OR = '0') then
         s_Energy_Bin_525 <= s_Energy_Bin_525 +'1';
		 Energy_Bin_Rdy_525 <= '1';
		else
		 s_Energy_Bin_525 <= s_Energy_Bin_525;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_525 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_525;  
 
  
  Energy_Bin_526 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_526   <=  (others =>'0');
		Energy_Bin_Rdy_526 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E526_C1_L and PEAK_C1 <= s_E526_C1_H and Bin_OR = '0') then
         s_Energy_Bin_526 <= s_Energy_Bin_526 +'1';
		 Energy_Bin_Rdy_526 <= '1';
		else
		 s_Energy_Bin_526 <= s_Energy_Bin_526;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_526 <= '0';
      end if;
    end if;
  end process  Energy_Bin_526;   
  
 Energy_Bin_527 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_527   <=  (others =>'0');
		Energy_Bin_Rdy_527 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E527_C1_L and PEAK_C1 <= s_E527_C1_H and Bin_OR = '0') then
         s_Energy_Bin_527 <= s_Energy_Bin_527 +'1';
		 Energy_Bin_Rdy_527 <= '1';
		else
		 s_Energy_Bin_527 <= s_Energy_Bin_527;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_527 <= '0';
      end if;
    end if;
  end process  Energy_Bin_527;   
  
  Energy_Bin_528 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_528   <=  (others =>'0');
		Energy_Bin_Rdy_528 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E528_C1_L and PEAK_C1 <= s_E528_C1_H and Bin_OR = '0') then
         s_Energy_Bin_528 <= s_Energy_Bin_528 +'1';
		 Energy_Bin_Rdy_528 <= '1';
		else
		 s_Energy_Bin_528 <= s_Energy_Bin_528;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_528 <= '0';
      end if;
    end if;
  end process  Energy_Bin_528;   
  
  Energy_Bin_529 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_529   <=  (others =>'0');
		Energy_Bin_Rdy_529 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E529_C1_L and PEAK_C1 <= s_E529_C1_H and Bin_OR = '0') then
         s_Energy_Bin_529 <= s_Energy_Bin_529 +'1';
		 Energy_Bin_Rdy_529 <= '1';
		else
		 s_Energy_Bin_529 <= s_Energy_Bin_529;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_529 <= '0';
      end if;
    end if;
  end process  Energy_Bin_529;        
  
     Energy_Bin_530 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_530   <=  (others =>'0');
		Energy_Bin_Rdy_530 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E530_C1_L and PEAK_C1 <= s_E530_C1_H and Bin_OR = '0') then
         s_Energy_Bin_530 <= s_Energy_Bin_530 +'1';
		 Energy_Bin_Rdy_530 <= '1';
		else
		 s_Energy_Bin_530 <= s_Energy_Bin_530;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_530 <= '0';
      end if;
    end if;
  end process  Energy_Bin_530;    
  
  Energy_Bin_531 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_531   <=  (others =>'0');
		Energy_Bin_Rdy_531 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E531_C1_L and PEAK_C1 <= s_E531_C1_H and Bin_OR = '0') then
         s_Energy_Bin_531 <= s_Energy_Bin_531 +'1';
		 Energy_Bin_Rdy_531 <= '1';
		else
		 s_Energy_Bin_531 <= s_Energy_Bin_531;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_531 <= '0';
      end if;
    end if;
  end process  Energy_Bin_531;   
  
  Energy_Bin_532 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_532   <=  (others =>'0');
	    Energy_Bin_Rdy_532 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E532_C1_L and PEAK_C1 <= s_E532_C1_H and Bin_OR = '0') then
         s_Energy_Bin_532 <= s_Energy_Bin_532 +'1';
		 Energy_Bin_Rdy_532 <= '1';
		else
		 s_Energy_Bin_532 <= s_Energy_Bin_532;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_532 <= '0';
      end if;
    end if;
  end process  Energy_Bin_532;   
  
  Energy_Bin_533 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_533   <=  (others =>'0');
	    Energy_Bin_Rdy_533 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E533_C1_L and PEAK_C1 <= s_E533_C1_H and Bin_OR = '0') then
         s_Energy_Bin_533 <= s_Energy_Bin_533 +'1';
		 Energy_Bin_Rdy_533 <= '1';
		else
		 s_Energy_Bin_533 <= s_Energy_Bin_533;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_533 <= '0';
      end if;
    end if;
  end process  Energy_Bin_533;   
  
  Energy_Bin_534 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_534   <=  (others =>'0');
		Energy_Bin_Rdy_534 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E534_C1_L and PEAK_C1 <= s_E534_C1_H and Bin_OR = '0') then
         s_Energy_Bin_534 <= s_Energy_Bin_534 +'1';
		 Energy_Bin_Rdy_534 <= '1';
		else
		 s_Energy_Bin_534 <= s_Energy_Bin_534;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_534 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_534;   
 
 
  Energy_Bin_535 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_535   <=  (others =>'0');
		Energy_Bin_Rdy_535 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E535_C1_L and PEAK_C1 <= s_E535_C1_H and Bin_OR = '0') then
         s_Energy_Bin_535 <= s_Energy_Bin_535 +'1';
		 Energy_Bin_Rdy_535 <= '1';
		else
		 s_Energy_Bin_535 <= s_Energy_Bin_535;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_535 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_535;  
 
  
  Energy_Bin_536 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_536   <=  (others =>'0');
		Energy_Bin_Rdy_536 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E536_C1_L and PEAK_C1 <= s_E536_C1_H and Bin_OR = '0') then
         s_Energy_Bin_536 <= s_Energy_Bin_536 +'1';
		 Energy_Bin_Rdy_536 <= '1';
		else
		 s_Energy_Bin_536 <= s_Energy_Bin_536;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_536 <= '0';
      end if;
    end if;
  end process  Energy_Bin_536;   
  
 Energy_Bin_537 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_537   <=  (others =>'0');
		Energy_Bin_Rdy_537 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E537_C1_L and PEAK_C1 <= s_E537_C1_H and Bin_OR = '0') then
         s_Energy_Bin_537 <= s_Energy_Bin_537 +'1';
		 Energy_Bin_Rdy_537 <= '1';
		else
		 s_Energy_Bin_537 <= s_Energy_Bin_537;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_537 <= '0';
      end if;
    end if;
  end process  Energy_Bin_537;   
  
  Energy_Bin_538 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_538   <=  (others =>'0');
		Energy_Bin_Rdy_538 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E538_C1_L and PEAK_C1 <= s_E538_C1_H and Bin_OR = '0') then
         s_Energy_Bin_538 <= s_Energy_Bin_538 +'1';
		 Energy_Bin_Rdy_538 <= '1';
		else
		 s_Energy_Bin_538 <= s_Energy_Bin_538;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_538 <= '0';
      end if;
    end if;
  end process  Energy_Bin_538;   
  
  Energy_Bin_539 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_539   <=  (others =>'0');
		Energy_Bin_Rdy_539 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E539_C1_L and PEAK_C1 <= s_E539_C1_H and Bin_OR = '0') then
         s_Energy_Bin_539 <= s_Energy_Bin_539 +'1';
		 Energy_Bin_Rdy_539 <= '1';
		else
		 s_Energy_Bin_539 <= s_Energy_Bin_539;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_539 <= '0';
      end if;
    end if;
  end process  Energy_Bin_539;         
  
     Energy_Bin_540 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_540   <=  (others =>'0');
		Energy_Bin_Rdy_540 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E540_C1_L and PEAK_C1 <= s_E540_C1_H and Bin_OR = '0') then
         s_Energy_Bin_540 <= s_Energy_Bin_540 +'1';
		 Energy_Bin_Rdy_540 <= '1';
		else
		 s_Energy_Bin_540 <= s_Energy_Bin_540;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_540 <= '0';
      end if;
    end if;
  end process  Energy_Bin_540;    
  
  Energy_Bin_541 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_541   <=  (others =>'0');
		Energy_Bin_Rdy_541 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E541_C1_L and PEAK_C1 <= s_E541_C1_H and Bin_OR = '0') then
         s_Energy_Bin_541 <= s_Energy_Bin_541 +'1';
		 Energy_Bin_Rdy_541 <= '1';
		else
		 s_Energy_Bin_541 <= s_Energy_Bin_541;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_541 <= '0';
      end if;
    end if;
  end process  Energy_Bin_541;   
  
  Energy_Bin_542 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_542   <=  (others =>'0');
	    Energy_Bin_Rdy_542 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E542_C1_L and PEAK_C1 <= s_E542_C1_H and Bin_OR = '0') then
         s_Energy_Bin_542 <= s_Energy_Bin_542 +'1';
		 Energy_Bin_Rdy_542 <= '1';
		else
		 s_Energy_Bin_542 <= s_Energy_Bin_542;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_542 <= '0';
      end if;
    end if;
  end process  Energy_Bin_542;   
  
  Energy_Bin_543 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_543   <=  (others =>'0');
	    Energy_Bin_Rdy_543 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E543_C1_L and PEAK_C1 <= s_E543_C1_H and Bin_OR = '0') then
         s_Energy_Bin_543 <= s_Energy_Bin_543 +'1';
		 Energy_Bin_Rdy_543 <= '1';
		else
		 s_Energy_Bin_543 <= s_Energy_Bin_543;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_543 <= '0';
      end if;
    end if;
  end process  Energy_Bin_543;   
  
  Energy_Bin_544 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_544   <=  (others =>'0');
		Energy_Bin_Rdy_544 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E544_C1_L and PEAK_C1 <= s_E544_C1_H and Bin_OR = '0') then
         s_Energy_Bin_544 <= s_Energy_Bin_544 +'1';
		 Energy_Bin_Rdy_544 <= '1';
		else
		 s_Energy_Bin_544 <= s_Energy_Bin_544;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_544 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_544;   
 
 
  Energy_Bin_545 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_545   <=  (others =>'0');
		Energy_Bin_Rdy_545 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E545_C1_L and PEAK_C1 <= s_E545_C1_H and Bin_OR = '0') then
         s_Energy_Bin_545 <= s_Energy_Bin_545 +'1';
		 Energy_Bin_Rdy_545 <= '1';
		else
		 s_Energy_Bin_545 <= s_Energy_Bin_545;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_545 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_545;  
 
  
  Energy_Bin_546 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_546   <=  (others =>'0');
		Energy_Bin_Rdy_546 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E546_C1_L and PEAK_C1 <= s_E546_C1_H and Bin_OR = '0') then
         s_Energy_Bin_546 <= s_Energy_Bin_546 +'1';
		 Energy_Bin_Rdy_546 <= '1';
		else
		 s_Energy_Bin_546 <= s_Energy_Bin_546;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_546 <= '0';
      end if;
    end if;
  end process  Energy_Bin_546;   
  
 Energy_Bin_547 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_547   <=  (others =>'0');
		Energy_Bin_Rdy_547 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E547_C1_L and PEAK_C1 <= s_E547_C1_H and Bin_OR = '0') then
         s_Energy_Bin_547 <= s_Energy_Bin_547 +'1';
		 Energy_Bin_Rdy_547 <= '1';
		else
		 s_Energy_Bin_547 <= s_Energy_Bin_547;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_547 <= '0';
      end if;
    end if;
  end process  Energy_Bin_547;   
  
  Energy_Bin_548 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_548   <=  (others =>'0');
		Energy_Bin_Rdy_548 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E548_C1_L and PEAK_C1 <= s_E548_C1_H and Bin_OR = '0') then
         s_Energy_Bin_548 <= s_Energy_Bin_548 +'1';
		 Energy_Bin_Rdy_548 <= '1';
		else
		 s_Energy_Bin_548 <= s_Energy_Bin_548;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_548 <= '0';
      end if;
    end if;
  end process  Energy_Bin_548;   
  
  Energy_Bin_549 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_549   <=  (others =>'0');
		Energy_Bin_Rdy_549 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E549_C1_L and PEAK_C1 <= s_E549_C1_H and Bin_OR = '0') then
         s_Energy_Bin_549 <= s_Energy_Bin_549 +'1';
		 Energy_Bin_Rdy_549 <= '1';
		else
		 s_Energy_Bin_549 <= s_Energy_Bin_549;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_549 <= '0';
      end if;
    end if;
  end process  Energy_Bin_549;          
  
  
     Energy_Bin_550 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_550   <=  (others =>'0');
		Energy_Bin_Rdy_550 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E550_C1_L and PEAK_C1 <= s_E550_C1_H and Bin_OR = '0') then
         s_Energy_Bin_550 <= s_Energy_Bin_550 +'1';
		 Energy_Bin_Rdy_550 <= '1';
		else
		 s_Energy_Bin_550 <= s_Energy_Bin_550;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_550 <= '0';
      end if;
    end if;
  end process  Energy_Bin_550;    
  
  Energy_Bin_551 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_551   <=  (others =>'0');
		Energy_Bin_Rdy_551 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E551_C1_L and PEAK_C1 <= s_E551_C1_H and Bin_OR = '0') then
         s_Energy_Bin_551 <= s_Energy_Bin_551 +'1';
		 Energy_Bin_Rdy_551 <= '1';
		else
		 s_Energy_Bin_551 <= s_Energy_Bin_551;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_551 <= '0';
      end if;
    end if;
  end process  Energy_Bin_551;   
  
  Energy_Bin_552 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_552   <=  (others =>'0');
	    Energy_Bin_Rdy_552 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E552_C1_L and PEAK_C1 <= s_E552_C1_H and Bin_OR = '0') then
         s_Energy_Bin_552 <= s_Energy_Bin_552 +'1';
		 Energy_Bin_Rdy_552 <= '1';
		else
		 s_Energy_Bin_552 <= s_Energy_Bin_552;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_552 <= '0';
      end if;
    end if;
  end process  Energy_Bin_552;   
  
  Energy_Bin_553 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_553   <=  (others =>'0');
	    Energy_Bin_Rdy_553 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E553_C1_L and PEAK_C1 <= s_E553_C1_H and Bin_OR = '0') then
         s_Energy_Bin_553 <= s_Energy_Bin_553 +'1';
		 Energy_Bin_Rdy_553 <= '1';
		else
		 s_Energy_Bin_553 <= s_Energy_Bin_553;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_553 <= '0';
      end if;
    end if;
  end process  Energy_Bin_553;   
  
  Energy_Bin_554 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_554   <=  (others =>'0');
		Energy_Bin_Rdy_554 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E554_C1_L and PEAK_C1 <= s_E554_C1_H and Bin_OR = '0') then
         s_Energy_Bin_554 <= s_Energy_Bin_554 +'1';
		 Energy_Bin_Rdy_554 <= '1';
		else
		 s_Energy_Bin_554 <= s_Energy_Bin_554;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_554 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_554;   
 
 
  Energy_Bin_555 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_555   <=  (others =>'0');
		Energy_Bin_Rdy_555 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E555_C1_L and PEAK_C1 <= s_E555_C1_H and Bin_OR = '0') then
         s_Energy_Bin_555 <= s_Energy_Bin_555 +'1';
		 Energy_Bin_Rdy_555 <= '1';
		else
		 s_Energy_Bin_555 <= s_Energy_Bin_555;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_555 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_555;  
 
  
  Energy_Bin_556 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_556   <=  (others =>'0');
		Energy_Bin_Rdy_556 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E556_C1_L and PEAK_C1 <= s_E556_C1_H and Bin_OR = '0') then
         s_Energy_Bin_556 <= s_Energy_Bin_556 +'1';
		 Energy_Bin_Rdy_556 <= '1';
		else
		 s_Energy_Bin_556 <= s_Energy_Bin_556;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_556 <= '0';
      end if;
    end if;
  end process  Energy_Bin_556;   
  
 Energy_Bin_557 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_557   <=  (others =>'0');
		Energy_Bin_Rdy_557 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E557_C1_L and PEAK_C1 <= s_E557_C1_H and Bin_OR = '0') then
         s_Energy_Bin_557 <= s_Energy_Bin_557 +'1';
		 Energy_Bin_Rdy_557 <= '1';
		else
		 s_Energy_Bin_557 <= s_Energy_Bin_557;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_557 <= '0';
      end if;
    end if;
  end process  Energy_Bin_557;   
  
  Energy_Bin_558 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_558   <=  (others =>'0');
		Energy_Bin_Rdy_558 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E558_C1_L and PEAK_C1 <= s_E558_C1_H and Bin_OR = '0') then
         s_Energy_Bin_558 <= s_Energy_Bin_558 +'1';
		 Energy_Bin_Rdy_558 <= '1';
		else
		 s_Energy_Bin_558 <= s_Energy_Bin_558;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_558 <= '0';
      end if;
    end if;
  end process  Energy_Bin_558;   
  
  Energy_Bin_559 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_559   <=  (others =>'0');
		Energy_Bin_Rdy_559 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E559_C1_L and PEAK_C1 <= s_E559_C1_H and Bin_OR = '0') then
         s_Energy_Bin_559 <= s_Energy_Bin_559 +'1';
		 Energy_Bin_Rdy_559 <= '1';
		else
		 s_Energy_Bin_559 <= s_Energy_Bin_559;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_559 <= '0';
      end if;
    end if;
  end process  Energy_Bin_559;           
  
     Energy_Bin_560 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_560   <=  (others =>'0');
		Energy_Bin_Rdy_560 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E560_C1_L and PEAK_C1 <= s_E560_C1_H and Bin_OR = '0') then
         s_Energy_Bin_560 <= s_Energy_Bin_560 +'1';
		 Energy_Bin_Rdy_560 <= '1';
		else
		 s_Energy_Bin_560 <= s_Energy_Bin_560;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_560 <= '0';
      end if;
    end if;
  end process  Energy_Bin_560;    
  
  Energy_Bin_561 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_561   <=  (others =>'0');
		Energy_Bin_Rdy_561 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E561_C1_L and PEAK_C1 <= s_E561_C1_H and Bin_OR = '0') then
         s_Energy_Bin_561 <= s_Energy_Bin_561 +'1';
		 Energy_Bin_Rdy_561 <= '1';
		else
		 s_Energy_Bin_561 <= s_Energy_Bin_561;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_561 <= '0';
      end if;
    end if;
  end process  Energy_Bin_561;   
  
  Energy_Bin_562 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_562   <=  (others =>'0');
	    Energy_Bin_Rdy_562 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E562_C1_L and PEAK_C1 <= s_E562_C1_H and Bin_OR = '0') then
         s_Energy_Bin_562 <= s_Energy_Bin_562 +'1';
		 Energy_Bin_Rdy_562 <= '1';
		else
		 s_Energy_Bin_562 <= s_Energy_Bin_562;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_562 <= '0';
      end if;
    end if;
  end process  Energy_Bin_562;   
  
  Energy_Bin_563 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_563   <=  (others =>'0');
	    Energy_Bin_Rdy_563 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E563_C1_L and PEAK_C1 <= s_E563_C1_H and Bin_OR = '0') then
         s_Energy_Bin_563 <= s_Energy_Bin_563 +'1';
		 Energy_Bin_Rdy_563 <= '1';
		else
		 s_Energy_Bin_563 <= s_Energy_Bin_563;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_563 <= '0';
      end if;
    end if;
  end process  Energy_Bin_563;   
  
  Energy_Bin_564 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_564   <=  (others =>'0');
		Energy_Bin_Rdy_564 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E564_C1_L and PEAK_C1 <= s_E564_C1_H and Bin_OR = '0') then
         s_Energy_Bin_564 <= s_Energy_Bin_564 +'1';
		 Energy_Bin_Rdy_564 <= '1';
		else
		 s_Energy_Bin_564 <= s_Energy_Bin_564;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_564 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_564;   
 
 
  Energy_Bin_565 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_565   <=  (others =>'0');
		Energy_Bin_Rdy_565 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E565_C1_L and PEAK_C1 <= s_E565_C1_H and Bin_OR = '0') then
         s_Energy_Bin_565 <= s_Energy_Bin_565 +'1';
		 Energy_Bin_Rdy_565 <= '1';
		else
		 s_Energy_Bin_565 <= s_Energy_Bin_565;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_565 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_565;  
 
  
  Energy_Bin_566 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_566   <=  (others =>'0');
		Energy_Bin_Rdy_566 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E566_C1_L and PEAK_C1 <= s_E566_C1_H and Bin_OR = '0') then
         s_Energy_Bin_566 <= s_Energy_Bin_566 +'1';
		 Energy_Bin_Rdy_566 <= '1';
		else
		 s_Energy_Bin_566 <= s_Energy_Bin_566;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_566 <= '0';
      end if;
    end if;
  end process  Energy_Bin_566;   
  
 Energy_Bin_567 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_567   <=  (others =>'0');
		Energy_Bin_Rdy_567 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E567_C1_L and PEAK_C1 <= s_E567_C1_H and Bin_OR = '0') then
         s_Energy_Bin_567 <= s_Energy_Bin_567 +'1';
		 Energy_Bin_Rdy_567 <= '1';
		else
		 s_Energy_Bin_567 <= s_Energy_Bin_567;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_567 <= '0';
      end if;
    end if;
  end process  Energy_Bin_567;   
  
  Energy_Bin_568 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_568   <=  (others =>'0');
		Energy_Bin_Rdy_568 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E568_C1_L and PEAK_C1 <= s_E568_C1_H and Bin_OR = '0') then
         s_Energy_Bin_568 <= s_Energy_Bin_568 +'1';
		 Energy_Bin_Rdy_568 <= '1';
		else
		 s_Energy_Bin_568 <= s_Energy_Bin_568;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_568 <= '0';
      end if;
    end if;
  end process  Energy_Bin_568;   
  
  Energy_Bin_569 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_569   <=  (others =>'0');
		Energy_Bin_Rdy_569 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E569_C1_L and PEAK_C1 <= s_E569_C1_H and Bin_OR = '0') then
         s_Energy_Bin_569 <= s_Energy_Bin_569 +'1';
		 Energy_Bin_Rdy_569 <= '1';
		else
		 s_Energy_Bin_569 <= s_Energy_Bin_569;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_569 <= '0';
      end if;
    end if;
  end process  Energy_Bin_569;         
  
     Energy_Bin_570 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_570   <=  (others =>'0');
		Energy_Bin_Rdy_570 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E570_C1_L and PEAK_C1 <= s_E570_C1_H and Bin_OR = '0') then
         s_Energy_Bin_570 <= s_Energy_Bin_570 +'1';
		 Energy_Bin_Rdy_570 <= '1';
		else
		 s_Energy_Bin_570 <= s_Energy_Bin_570;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_570 <= '0';
      end if;
    end if;
  end process  Energy_Bin_570;    
  
  Energy_Bin_571 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_571   <=  (others =>'0');
		Energy_Bin_Rdy_571 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E571_C1_L and PEAK_C1 <= s_E571_C1_H and Bin_OR = '0') then
         s_Energy_Bin_571 <= s_Energy_Bin_571 +'1';
		 Energy_Bin_Rdy_571 <= '1';
		else
		 s_Energy_Bin_571 <= s_Energy_Bin_571;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_571 <= '0';
      end if;
    end if;
  end process  Energy_Bin_571;   
  
  Energy_Bin_572 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_572   <=  (others =>'0');
	    Energy_Bin_Rdy_572 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E572_C1_L and PEAK_C1 <= s_E572_C1_H and Bin_OR = '0') then
         s_Energy_Bin_572 <= s_Energy_Bin_572 +'1';
		 Energy_Bin_Rdy_572 <= '1';
		else
		 s_Energy_Bin_572 <= s_Energy_Bin_572;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_572 <= '0';
      end if;
    end if;
  end process  Energy_Bin_572;   
  
  Energy_Bin_573 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_573   <=  (others =>'0');
	    Energy_Bin_Rdy_573 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E573_C1_L and PEAK_C1 <= s_E573_C1_H and Bin_OR = '0') then
         s_Energy_Bin_573 <= s_Energy_Bin_573 +'1';
		 Energy_Bin_Rdy_573 <= '1';
		else
		 s_Energy_Bin_573 <= s_Energy_Bin_573;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_573 <= '0';
      end if;
    end if;
  end process  Energy_Bin_573;   
  
  Energy_Bin_574 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_574   <=  (others =>'0');
		Energy_Bin_Rdy_574 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E574_C1_L and PEAK_C1 <= s_E574_C1_H and Bin_OR = '0') then
         s_Energy_Bin_574 <= s_Energy_Bin_574 +'1';
		 Energy_Bin_Rdy_574 <= '1';
		else
		 s_Energy_Bin_574 <= s_Energy_Bin_574;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_574 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_574;   
 
 
  Energy_Bin_575 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_575   <=  (others =>'0');
		Energy_Bin_Rdy_575 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E575_C1_L and PEAK_C1 <= s_E575_C1_H and Bin_OR = '0') then
         s_Energy_Bin_575 <= s_Energy_Bin_575 +'1';
		 Energy_Bin_Rdy_575 <= '1';
		else
		 s_Energy_Bin_575 <= s_Energy_Bin_575;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_575 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_575;  
 
  
  Energy_Bin_576 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_576   <=  (others =>'0');
		Energy_Bin_Rdy_576 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E576_C1_L and PEAK_C1 <= s_E576_C1_H and Bin_OR = '0') then
         s_Energy_Bin_576 <= s_Energy_Bin_576 +'1';
		 Energy_Bin_Rdy_576 <= '1';
		else
		 s_Energy_Bin_576 <= s_Energy_Bin_576;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_576 <= '0';
      end if;
    end if;
  end process  Energy_Bin_576;   
  
 Energy_Bin_577 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_577   <=  (others =>'0');
		Energy_Bin_Rdy_577 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E577_C1_L and PEAK_C1 <= s_E577_C1_H and Bin_OR = '0') then
         s_Energy_Bin_577 <= s_Energy_Bin_577 +'1';
		 Energy_Bin_Rdy_577 <= '1';
		else
		 s_Energy_Bin_577 <= s_Energy_Bin_577;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_577 <= '0';
      end if;
    end if;
  end process  Energy_Bin_577;   
  
  Energy_Bin_578 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_578   <=  (others =>'0');
		Energy_Bin_Rdy_578 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E578_C1_L and PEAK_C1 <= s_E578_C1_H and Bin_OR = '0') then
         s_Energy_Bin_578 <= s_Energy_Bin_578 +'1';
		 Energy_Bin_Rdy_578 <= '1';
		else
		 s_Energy_Bin_578 <= s_Energy_Bin_578;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_578 <= '0';
      end if;
    end if;
  end process  Energy_Bin_578;   
  
  Energy_Bin_579 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_579   <=  (others =>'0');
		Energy_Bin_Rdy_579 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E579_C1_L and PEAK_C1 <= s_E579_C1_H and Bin_OR = '0') then
         s_Energy_Bin_579 <= s_Energy_Bin_579 +'1';
		 Energy_Bin_Rdy_579 <= '1';
		else
		 s_Energy_Bin_579 <= s_Energy_Bin_579;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_579 <= '0';
      end if;
    end if;
  end process  Energy_Bin_579;       
  
     Energy_Bin_580 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_580   <=  (others =>'0');
		Energy_Bin_Rdy_580 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E580_C1_L and PEAK_C1 <= s_E580_C1_H and Bin_OR = '0') then
         s_Energy_Bin_580 <= s_Energy_Bin_580 +'1';
		 Energy_Bin_Rdy_580 <= '1';
		else
		 s_Energy_Bin_580 <= s_Energy_Bin_580;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_580 <= '0';
      end if;
    end if;
  end process  Energy_Bin_580;    
  
  Energy_Bin_581 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_581   <=  (others =>'0');
		Energy_Bin_Rdy_581 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E581_C1_L and PEAK_C1 <= s_E581_C1_H and Bin_OR = '0') then
         s_Energy_Bin_581 <= s_Energy_Bin_581 +'1';
		 Energy_Bin_Rdy_581 <= '1';
		else
		 s_Energy_Bin_581 <= s_Energy_Bin_581;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_581 <= '0';
      end if;
    end if;
  end process  Energy_Bin_581;   
  
  Energy_Bin_582 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_582   <=  (others =>'0');
	    Energy_Bin_Rdy_582 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E582_C1_L and PEAK_C1 <= s_E582_C1_H and Bin_OR = '0') then
         s_Energy_Bin_582 <= s_Energy_Bin_582 +'1';
		 Energy_Bin_Rdy_582 <= '1';
		else
		 s_Energy_Bin_582 <= s_Energy_Bin_582;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_582 <= '0';
      end if;
    end if;
  end process  Energy_Bin_582;   
  
  Energy_Bin_583 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_583   <=  (others =>'0');
	    Energy_Bin_Rdy_583 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E583_C1_L and PEAK_C1 <= s_E583_C1_H and Bin_OR = '0') then
         s_Energy_Bin_583 <= s_Energy_Bin_583 +'1';
		 Energy_Bin_Rdy_583 <= '1';
		else
		 s_Energy_Bin_583 <= s_Energy_Bin_583;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_583 <= '0';
      end if;
    end if;
  end process  Energy_Bin_583;   
  
  Energy_Bin_584 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_584   <=  (others =>'0');
		Energy_Bin_Rdy_584 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E584_C1_L and PEAK_C1 <= s_E584_C1_H and Bin_OR = '0') then
         s_Energy_Bin_584 <= s_Energy_Bin_584 +'1';
		 Energy_Bin_Rdy_584 <= '1';
		else
		 s_Energy_Bin_584 <= s_Energy_Bin_584;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_584 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_584;   
 
 
  Energy_Bin_585 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_585   <=  (others =>'0');
		Energy_Bin_Rdy_585 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E585_C1_L and PEAK_C1 <= s_E585_C1_H and Bin_OR = '0') then
         s_Energy_Bin_585 <= s_Energy_Bin_585 +'1';
		 Energy_Bin_Rdy_585 <= '1';
		else
		 s_Energy_Bin_585 <= s_Energy_Bin_585;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_585 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_585;  
 
  
  Energy_Bin_586 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_586   <=  (others =>'0');
		Energy_Bin_Rdy_586 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E586_C1_L and PEAK_C1 <= s_E586_C1_H and Bin_OR = '0') then
         s_Energy_Bin_586 <= s_Energy_Bin_586 +'1';
		 Energy_Bin_Rdy_586 <= '1';
		else
		 s_Energy_Bin_586 <= s_Energy_Bin_586;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_586 <= '0';
      end if;
    end if;
  end process  Energy_Bin_586;   
  
 Energy_Bin_587 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_587   <=  (others =>'0');
		Energy_Bin_Rdy_587 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E587_C1_L and PEAK_C1 <= s_E587_C1_H and Bin_OR = '0') then
         s_Energy_Bin_587 <= s_Energy_Bin_587 +'1';
		 Energy_Bin_Rdy_587 <= '1';
		else
		 s_Energy_Bin_587 <= s_Energy_Bin_587;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_587 <= '0';
      end if;
    end if;
  end process  Energy_Bin_587;   
  
  Energy_Bin_588 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_588   <=  (others =>'0');
		Energy_Bin_Rdy_588 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E588_C1_L and PEAK_C1 <= s_E588_C1_H and Bin_OR = '0') then
         s_Energy_Bin_588 <= s_Energy_Bin_588 +'1';
		 Energy_Bin_Rdy_588 <= '1';
		else
		 s_Energy_Bin_588 <= s_Energy_Bin_588;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_588 <= '0';
      end if;
    end if;
  end process  Energy_Bin_588;   
  
  Energy_Bin_589 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_589   <=  (others =>'0');
		Energy_Bin_Rdy_589 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E589_C1_L and PEAK_C1 <= s_E589_C1_H and Bin_OR = '0') then
         s_Energy_Bin_589 <= s_Energy_Bin_589 +'1';
		 Energy_Bin_Rdy_589 <= '1';
		else
		 s_Energy_Bin_589 <= s_Energy_Bin_589;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_589 <= '0';
      end if;
    end if;
  end process  Energy_Bin_589;      
  
     Energy_Bin_590 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_590   <=  (others =>'0');
		Energy_Bin_Rdy_590 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E590_C1_L and PEAK_C1 <= s_E590_C1_H and Bin_OR = '0') then
         s_Energy_Bin_590 <= s_Energy_Bin_590 +'1';
		 Energy_Bin_Rdy_590 <= '1';
		else
		 s_Energy_Bin_590 <= s_Energy_Bin_590;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_590 <= '0';
      end if;
    end if;
  end process  Energy_Bin_590;    
  
  Energy_Bin_591 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_591   <=  (others =>'0');
		Energy_Bin_Rdy_591 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E591_C1_L and PEAK_C1 <= s_E591_C1_H and Bin_OR = '0') then
         s_Energy_Bin_591 <= s_Energy_Bin_591 +'1';
		 Energy_Bin_Rdy_591 <= '1';
		else
		 s_Energy_Bin_591 <= s_Energy_Bin_591;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_591 <= '0';
      end if;
    end if;
  end process  Energy_Bin_591;   
  
  Energy_Bin_592 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_592   <=  (others =>'0');
	    Energy_Bin_Rdy_592 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E592_C1_L and PEAK_C1 <= s_E592_C1_H and Bin_OR = '0') then
         s_Energy_Bin_592 <= s_Energy_Bin_592 +'1';
		 Energy_Bin_Rdy_592 <= '1';
		else
		 s_Energy_Bin_592 <= s_Energy_Bin_592;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_592 <= '0';
      end if;
    end if;
  end process  Energy_Bin_592;   
  
  Energy_Bin_593 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_593   <=  (others =>'0');
	    Energy_Bin_Rdy_593 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E593_C1_L and PEAK_C1 <= s_E593_C1_H and Bin_OR = '0') then
         s_Energy_Bin_593 <= s_Energy_Bin_593 +'1';
		 Energy_Bin_Rdy_593 <= '1';
		else
		 s_Energy_Bin_593 <= s_Energy_Bin_593;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_593 <= '0';
      end if;
    end if;
  end process  Energy_Bin_593;   
  
  Energy_Bin_594 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_594   <=  (others =>'0');
		Energy_Bin_Rdy_594 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E594_C1_L and PEAK_C1 <= s_E594_C1_H and Bin_OR = '0') then
         s_Energy_Bin_594 <= s_Energy_Bin_594 +'1';
		 Energy_Bin_Rdy_594 <= '1';
		else
		 s_Energy_Bin_594 <= s_Energy_Bin_594;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_594 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_594;   
 
 
  Energy_Bin_595 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_595   <=  (others =>'0');
		Energy_Bin_Rdy_595 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E595_C1_L and PEAK_C1 <= s_E595_C1_H and Bin_OR = '0') then
         s_Energy_Bin_595 <= s_Energy_Bin_595 +'1';
		 Energy_Bin_Rdy_595 <= '1';
		else
		 s_Energy_Bin_595 <= s_Energy_Bin_595;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_595 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_595;  
 
  
  Energy_Bin_596 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_596   <=  (others =>'0');
		Energy_Bin_Rdy_596 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E596_C1_L and PEAK_C1 <= s_E596_C1_H and Bin_OR = '0') then
         s_Energy_Bin_596 <= s_Energy_Bin_596 +'1';
		 Energy_Bin_Rdy_596 <= '1';
		else
		 s_Energy_Bin_596 <= s_Energy_Bin_596;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_596 <= '0';
      end if;
    end if;
  end process  Energy_Bin_596;   
  
 Energy_Bin_597 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_597   <=  (others =>'0');
		Energy_Bin_Rdy_597 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E597_C1_L and PEAK_C1 <= s_E597_C1_H and Bin_OR = '0') then
         s_Energy_Bin_597 <= s_Energy_Bin_597 +'1';
		 Energy_Bin_Rdy_597 <= '1';
		else
		 s_Energy_Bin_597 <= s_Energy_Bin_597;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_597 <= '0';
      end if;
    end if;
  end process  Energy_Bin_597;   
  
  Energy_Bin_598 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_598   <=  (others =>'0');
		Energy_Bin_Rdy_598 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E598_C1_L and PEAK_C1 <= s_E598_C1_H and Bin_OR = '0') then
         s_Energy_Bin_598 <= s_Energy_Bin_598 +'1';
		 Energy_Bin_Rdy_598 <= '1';
		else
		 s_Energy_Bin_598 <= s_Energy_Bin_598;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_598 <= '0';
      end if;
    end if;
  end process  Energy_Bin_598;   
  
  Energy_Bin_599 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_599   <=  (others =>'0');
		Energy_Bin_Rdy_599 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E599_C1_L and PEAK_C1 <= s_E599_C1_H and Bin_OR = '0') then
         s_Energy_Bin_599 <= s_Energy_Bin_599 +'1';
		 Energy_Bin_Rdy_599 <= '1';
		else
		 s_Energy_Bin_599 <= s_Energy_Bin_599;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_599 <= '0';
      end if;
    end if;
  end process  Energy_Bin_599;      

    Energy_Bin_600 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_600   <=  (others =>'0');
		Energy_Bin_Rdy_600 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E600_C1_L and PEAK_C1 <= s_E600_C1_H and Bin_OR = '0') then
         s_Energy_Bin_600 <= s_Energy_Bin_600 +'1';
		 Energy_Bin_Rdy_600 <= '1';
		else
		 s_Energy_Bin_600 <= s_Energy_Bin_600;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_600 <= '0';
      end if;
    end if;
  end process  Energy_Bin_600;    
  
  Energy_Bin_601 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_601   <=  (others =>'0');
		Energy_Bin_Rdy_601 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E601_C1_L and PEAK_C1 <= s_E601_C1_H and Bin_OR = '0') then
         s_Energy_Bin_601 <= s_Energy_Bin_601 +'1';
		 Energy_Bin_Rdy_601 <= '1';
		else
		 s_Energy_Bin_601 <= s_Energy_Bin_601;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_601 <= '0';
      end if;
    end if;
  end process  Energy_Bin_601;   
  
  Energy_Bin_602 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_602   <=  (others =>'0');
	    Energy_Bin_Rdy_602 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E602_C1_L and PEAK_C1 <= s_E602_C1_H and Bin_OR = '0') then
         s_Energy_Bin_602 <= s_Energy_Bin_602 +'1';
		 Energy_Bin_Rdy_602 <= '1';
		else
		 s_Energy_Bin_602 <= s_Energy_Bin_602;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_602 <= '0';
      end if;
    end if;
  end process  Energy_Bin_602;   
  
  Energy_Bin_603 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_603   <=  (others =>'0');
	    Energy_Bin_Rdy_603 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E603_C1_L and PEAK_C1 <= s_E603_C1_H and Bin_OR = '0') then
         s_Energy_Bin_603 <= s_Energy_Bin_603 +'1';
		 Energy_Bin_Rdy_603 <= '1';
		else
		 s_Energy_Bin_603 <= s_Energy_Bin_603;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_603 <= '0';
      end if;
    end if;
  end process  Energy_Bin_603;   
  
  Energy_Bin_604 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_604   <=  (others =>'0');
		Energy_Bin_Rdy_604 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E604_C1_L and PEAK_C1 <= s_E604_C1_H and Bin_OR = '0') then
         s_Energy_Bin_604 <= s_Energy_Bin_604 +'1';
		 Energy_Bin_Rdy_604 <= '1';
		else
		 s_Energy_Bin_604 <= s_Energy_Bin_604;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_604 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_604;   
 
 
  Energy_Bin_605 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_605   <=  (others =>'0');
		Energy_Bin_Rdy_605 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E605_C1_L and PEAK_C1 <= s_E605_C1_H and Bin_OR = '0') then
         s_Energy_Bin_605 <= s_Energy_Bin_605 +'1';
		 Energy_Bin_Rdy_605 <= '1';
		else
		 s_Energy_Bin_605 <= s_Energy_Bin_605;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_605 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_605;  
 
  
  Energy_Bin_606 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_606   <=  (others =>'0');
		Energy_Bin_Rdy_606 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E606_C1_L and PEAK_C1 <= s_E606_C1_H and Bin_OR = '0') then
         s_Energy_Bin_606 <= s_Energy_Bin_606 +'1';
		 Energy_Bin_Rdy_606 <= '1';
		else
		 s_Energy_Bin_606 <= s_Energy_Bin_606;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_606 <= '0';
      end if;
    end if;
  end process  Energy_Bin_606;   
  
 Energy_Bin_607 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_607   <=  (others =>'0');
		Energy_Bin_Rdy_607 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E607_C1_L and PEAK_C1 <= s_E607_C1_H and Bin_OR = '0') then
         s_Energy_Bin_607 <= s_Energy_Bin_607 +'1';
		 Energy_Bin_Rdy_607 <= '1';
		else
		 s_Energy_Bin_607 <= s_Energy_Bin_607;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_607 <= '0';
      end if;
    end if;
  end process  Energy_Bin_607;   
  
  Energy_Bin_608 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_608   <=  (others =>'0');
		Energy_Bin_Rdy_608 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E608_C1_L and PEAK_C1 <= s_E608_C1_H and Bin_OR = '0') then
         s_Energy_Bin_608 <= s_Energy_Bin_608 +'1';
		 Energy_Bin_Rdy_608 <= '1';
		else
		 s_Energy_Bin_608 <= s_Energy_Bin_608;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_608 <= '0';
      end if;
    end if;
  end process  Energy_Bin_608;   
  
  Energy_Bin_609 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_609   <=  (others =>'0');
		Energy_Bin_Rdy_609 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E609_C1_L and PEAK_C1 <= s_E609_C1_H and Bin_OR = '0') then
         s_Energy_Bin_609 <= s_Energy_Bin_609 +'1';
		 Energy_Bin_Rdy_609 <= '1';
		else
		 s_Energy_Bin_609 <= s_Energy_Bin_609;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_609 <= '0';
      end if;
    end if;
  end process  Energy_Bin_609;      
  
     Energy_Bin_610 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_610   <=  (others =>'0');
		Energy_Bin_Rdy_610 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E610_C1_L and PEAK_C1 <= s_E610_C1_H and Bin_OR = '0') then
         s_Energy_Bin_610 <= s_Energy_Bin_610 +'1';
		 Energy_Bin_Rdy_610 <= '1';
		else
		 s_Energy_Bin_610 <= s_Energy_Bin_610;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_610 <= '0';
      end if;
    end if;
  end process  Energy_Bin_610;    
  
  Energy_Bin_611 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_611   <=  (others =>'0');
		Energy_Bin_Rdy_611 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E611_C1_L and PEAK_C1 <= s_E611_C1_H and Bin_OR = '0') then
         s_Energy_Bin_611 <= s_Energy_Bin_611 +'1';
		 Energy_Bin_Rdy_611 <= '1';
		else
		 s_Energy_Bin_611 <= s_Energy_Bin_611;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_611 <= '0';
      end if;
    end if;
  end process  Energy_Bin_611;   
  
  Energy_Bin_612 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_612   <=  (others =>'0');
	    Energy_Bin_Rdy_612 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E612_C1_L and PEAK_C1 <= s_E612_C1_H and Bin_OR = '0') then
         s_Energy_Bin_612 <= s_Energy_Bin_612 +'1';
		 Energy_Bin_Rdy_612 <= '1';
		else
		 s_Energy_Bin_612 <= s_Energy_Bin_612;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_612 <= '0';
      end if;
    end if;
  end process  Energy_Bin_612;   
  
  Energy_Bin_613 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_613   <=  (others =>'0');
	    Energy_Bin_Rdy_613 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E613_C1_L and PEAK_C1 <= s_E613_C1_H and Bin_OR = '0') then
         s_Energy_Bin_613 <= s_Energy_Bin_613 +'1';
		 Energy_Bin_Rdy_613 <= '1';
		else
		 s_Energy_Bin_613 <= s_Energy_Bin_613;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_613 <= '0';
      end if;
    end if;
  end process  Energy_Bin_613;   
  
  Energy_Bin_614 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_614   <=  (others =>'0');
		Energy_Bin_Rdy_614 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E614_C1_L and PEAK_C1 <= s_E614_C1_H and Bin_OR = '0') then
         s_Energy_Bin_614 <= s_Energy_Bin_614 +'1';
		 Energy_Bin_Rdy_614 <= '1';
		else
		 s_Energy_Bin_614 <= s_Energy_Bin_614;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_614 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_614;   
 
 
  Energy_Bin_615 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_615   <=  (others =>'0');
		Energy_Bin_Rdy_615 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E615_C1_L and PEAK_C1 <= s_E615_C1_H and Bin_OR = '0') then
         s_Energy_Bin_615 <= s_Energy_Bin_615 +'1';
		 Energy_Bin_Rdy_615 <= '1';
		else
		 s_Energy_Bin_615 <= s_Energy_Bin_615;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_615 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_615;  
 
  
  Energy_Bin_616 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_616   <=  (others =>'0');
		Energy_Bin_Rdy_616 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E616_C1_L and PEAK_C1 <= s_E616_C1_H and Bin_OR = '0') then
         s_Energy_Bin_616 <= s_Energy_Bin_616 +'1';
		 Energy_Bin_Rdy_616 <= '1';
		else
		 s_Energy_Bin_616 <= s_Energy_Bin_616;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_616 <= '0';
      end if;
    end if;
  end process  Energy_Bin_616;   
  
 Energy_Bin_617 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_617   <=  (others =>'0');
		Energy_Bin_Rdy_617 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E617_C1_L and PEAK_C1 <= s_E617_C1_H and Bin_OR = '0') then
         s_Energy_Bin_617 <= s_Energy_Bin_617 +'1';
		 Energy_Bin_Rdy_617 <= '1';
		else
		 s_Energy_Bin_617 <= s_Energy_Bin_617;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_617 <= '0';
      end if;
    end if;
  end process  Energy_Bin_617;   
  
  Energy_Bin_618 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_618   <=  (others =>'0');
		Energy_Bin_Rdy_618 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E618_C1_L and PEAK_C1 <= s_E618_C1_H and Bin_OR = '0') then
         s_Energy_Bin_618 <= s_Energy_Bin_618 +'1';
		 Energy_Bin_Rdy_618 <= '1';
		else
		 s_Energy_Bin_618 <= s_Energy_Bin_618;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_618 <= '0';
      end if;
    end if;
  end process  Energy_Bin_618;   
  
  Energy_Bin_619 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_619   <=  (others =>'0');
		Energy_Bin_Rdy_619 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E619_C1_L and PEAK_C1 <= s_E619_C1_H and Bin_OR = '0') then
         s_Energy_Bin_619 <= s_Energy_Bin_619 +'1';
		 Energy_Bin_Rdy_619 <= '1';
		else
		 s_Energy_Bin_619 <= s_Energy_Bin_619;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_619 <= '0';
      end if;
    end if;
  end process  Energy_Bin_619;       
  
     Energy_Bin_620 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_620   <=  (others =>'0');
		Energy_Bin_Rdy_620 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E620_C1_L and PEAK_C1 <= s_E620_C1_H and Bin_OR = '0') then
         s_Energy_Bin_620 <= s_Energy_Bin_620 +'1';
		 Energy_Bin_Rdy_620 <= '1';
		else
		 s_Energy_Bin_620 <= s_Energy_Bin_620;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_620 <= '0';
      end if;
    end if;
  end process  Energy_Bin_620;    
  
  Energy_Bin_621 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_621   <=  (others =>'0');
		Energy_Bin_Rdy_621 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E621_C1_L and PEAK_C1 <= s_E621_C1_H and Bin_OR = '0') then
         s_Energy_Bin_621 <= s_Energy_Bin_621 +'1';
		 Energy_Bin_Rdy_621 <= '1';
		else
		 s_Energy_Bin_621 <= s_Energy_Bin_621;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_621 <= '0';
      end if;
    end if;
  end process  Energy_Bin_621;   
  
  Energy_Bin_622 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_622   <=  (others =>'0');
	    Energy_Bin_Rdy_622 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E622_C1_L and PEAK_C1 <= s_E622_C1_H and Bin_OR = '0') then
         s_Energy_Bin_622 <= s_Energy_Bin_622 +'1';
		 Energy_Bin_Rdy_622 <= '1';
		else
		 s_Energy_Bin_622 <= s_Energy_Bin_622;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_622 <= '0';
      end if;
    end if;
  end process  Energy_Bin_622;   
  
  Energy_Bin_623 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_623   <=  (others =>'0');
	    Energy_Bin_Rdy_623 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E623_C1_L and PEAK_C1 <= s_E623_C1_H and Bin_OR = '0') then
         s_Energy_Bin_623 <= s_Energy_Bin_623 +'1';
		 Energy_Bin_Rdy_623 <= '1';
		else
		 s_Energy_Bin_623 <= s_Energy_Bin_623;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_623 <= '0';
      end if;
    end if;
  end process  Energy_Bin_623;   
  
  Energy_Bin_624 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_624   <=  (others =>'0');
		Energy_Bin_Rdy_624 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E624_C1_L and PEAK_C1 <= s_E624_C1_H and Bin_OR = '0') then
         s_Energy_Bin_624 <= s_Energy_Bin_624 +'1';
		 Energy_Bin_Rdy_624 <= '1';
		else
		 s_Energy_Bin_624 <= s_Energy_Bin_624;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_624 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_624;   
 
 
  Energy_Bin_625 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_625   <=  (others =>'0');
		Energy_Bin_Rdy_625 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E625_C1_L and PEAK_C1 <= s_E625_C1_H and Bin_OR = '0') then
         s_Energy_Bin_625 <= s_Energy_Bin_625 +'1';
		 Energy_Bin_Rdy_625 <= '1';
		else
		 s_Energy_Bin_625 <= s_Energy_Bin_625;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_625 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_625;  
 
  
  Energy_Bin_626 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_626   <=  (others =>'0');
		Energy_Bin_Rdy_626 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E626_C1_L and PEAK_C1 <= s_E626_C1_H and Bin_OR = '0') then
         s_Energy_Bin_626 <= s_Energy_Bin_626 +'1';
		 Energy_Bin_Rdy_626 <= '1';
		else
		 s_Energy_Bin_626 <= s_Energy_Bin_626;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_626 <= '0';
      end if;
    end if;
  end process  Energy_Bin_626;   
  
 Energy_Bin_627 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_627   <=  (others =>'0');
		Energy_Bin_Rdy_627 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E627_C1_L and PEAK_C1 <= s_E627_C1_H and Bin_OR = '0') then
         s_Energy_Bin_627 <= s_Energy_Bin_627 +'1';
		 Energy_Bin_Rdy_627 <= '1';
		else
		 s_Energy_Bin_627 <= s_Energy_Bin_627;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_627 <= '0';
      end if;
    end if;
  end process  Energy_Bin_627;   
  
  Energy_Bin_628 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_628   <=  (others =>'0');
		Energy_Bin_Rdy_628 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E628_C1_L and PEAK_C1 <= s_E628_C1_H and Bin_OR = '0') then
         s_Energy_Bin_628 <= s_Energy_Bin_628 +'1';
		 Energy_Bin_Rdy_628 <= '1';
		else
		 s_Energy_Bin_628 <= s_Energy_Bin_628;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_628 <= '0';
      end if;
    end if;
  end process  Energy_Bin_628;   
  
  Energy_Bin_629 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_629   <=  (others =>'0');
		Energy_Bin_Rdy_629 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E629_C1_L and PEAK_C1 <= s_E629_C1_H and Bin_OR = '0') then
         s_Energy_Bin_629 <= s_Energy_Bin_629 +'1';
		 Energy_Bin_Rdy_629 <= '1';
		else
		 s_Energy_Bin_629 <= s_Energy_Bin_629;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_629 <= '0';
      end if;
    end if;
  end process  Energy_Bin_629;        
  
     Energy_Bin_630 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_630   <=  (others =>'0');
		Energy_Bin_Rdy_630 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E630_C1_L and PEAK_C1 <= s_E630_C1_H and Bin_OR = '0') then
         s_Energy_Bin_630 <= s_Energy_Bin_630 +'1';
		 Energy_Bin_Rdy_630 <= '1';
		else
		 s_Energy_Bin_630 <= s_Energy_Bin_630;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_630 <= '0';
      end if;
    end if;
  end process  Energy_Bin_630;    
  
  Energy_Bin_631 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_631   <=  (others =>'0');
		Energy_Bin_Rdy_631 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E631_C1_L and PEAK_C1 <= s_E631_C1_H and Bin_OR = '0') then
         s_Energy_Bin_631 <= s_Energy_Bin_631 +'1';
		 Energy_Bin_Rdy_631 <= '1';
		else
		 s_Energy_Bin_631 <= s_Energy_Bin_631;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_631 <= '0';
      end if;
    end if;
  end process  Energy_Bin_631;   
  
  Energy_Bin_632 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_632   <=  (others =>'0');
	    Energy_Bin_Rdy_632 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E632_C1_L and PEAK_C1 <= s_E632_C1_H and Bin_OR = '0') then
         s_Energy_Bin_632 <= s_Energy_Bin_632 +'1';
		 Energy_Bin_Rdy_632 <= '1';
		else
		 s_Energy_Bin_632 <= s_Energy_Bin_632;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_632 <= '0';
      end if;
    end if;
  end process  Energy_Bin_632;   
  
  Energy_Bin_633 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_633   <=  (others =>'0');
	    Energy_Bin_Rdy_633 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E633_C1_L and PEAK_C1 <= s_E633_C1_H and Bin_OR = '0') then
         s_Energy_Bin_633 <= s_Energy_Bin_633 +'1';
		 Energy_Bin_Rdy_633 <= '1';
		else
		 s_Energy_Bin_633 <= s_Energy_Bin_633;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_633 <= '0';
      end if;
    end if;
  end process  Energy_Bin_633;   
  
  Energy_Bin_634 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_634   <=  (others =>'0');
		Energy_Bin_Rdy_634 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E634_C1_L and PEAK_C1 <= s_E634_C1_H and Bin_OR = '0') then
         s_Energy_Bin_634 <= s_Energy_Bin_634 +'1';
		 Energy_Bin_Rdy_634 <= '1';
		else
		 s_Energy_Bin_634 <= s_Energy_Bin_634;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_634 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_634;   
 
 
  Energy_Bin_635 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_635   <=  (others =>'0');
		Energy_Bin_Rdy_635 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E635_C1_L and PEAK_C1 <= s_E635_C1_H and Bin_OR = '0') then
         s_Energy_Bin_635 <= s_Energy_Bin_635 +'1';
		 Energy_Bin_Rdy_635 <= '1';
		else
		 s_Energy_Bin_635 <= s_Energy_Bin_635;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_635 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_635;  
 
  
  Energy_Bin_636 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_636   <=  (others =>'0');
		Energy_Bin_Rdy_636 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E636_C1_L and PEAK_C1 <= s_E636_C1_H and Bin_OR = '0') then
         s_Energy_Bin_636 <= s_Energy_Bin_636 +'1';
		 Energy_Bin_Rdy_636 <= '1';
		else
		 s_Energy_Bin_636 <= s_Energy_Bin_636;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_636 <= '0';
      end if;
    end if;
  end process  Energy_Bin_636;   
  
 Energy_Bin_637 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_637   <=  (others =>'0');
		Energy_Bin_Rdy_637 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E637_C1_L and PEAK_C1 <= s_E637_C1_H and Bin_OR = '0') then
         s_Energy_Bin_637 <= s_Energy_Bin_637 +'1';
		 Energy_Bin_Rdy_637 <= '1';
		else
		 s_Energy_Bin_637 <= s_Energy_Bin_637;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_637 <= '0';
      end if;
    end if;
  end process  Energy_Bin_637;   
  
  Energy_Bin_638 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_638   <=  (others =>'0');
		Energy_Bin_Rdy_638 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E638_C1_L and PEAK_C1 <= s_E638_C1_H and Bin_OR = '0') then
         s_Energy_Bin_638 <= s_Energy_Bin_638 +'1';
		 Energy_Bin_Rdy_638 <= '1';
		else
		 s_Energy_Bin_638 <= s_Energy_Bin_638;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_638 <= '0';
      end if;
    end if;
  end process  Energy_Bin_638;   
  
  Energy_Bin_639 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_639   <=  (others =>'0');
		Energy_Bin_Rdy_639 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E639_C1_L and PEAK_C1 <= s_E639_C1_H and Bin_OR = '0') then
         s_Energy_Bin_639 <= s_Energy_Bin_639 +'1';
		 Energy_Bin_Rdy_639 <= '1';
		else
		 s_Energy_Bin_639 <= s_Energy_Bin_639;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_639 <= '0';
      end if;
    end if;
  end process  Energy_Bin_639;         
  
     Energy_Bin_640 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_640   <=  (others =>'0');
		Energy_Bin_Rdy_640 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E640_C1_L and PEAK_C1 <= s_E640_C1_H and Bin_OR = '0') then
         s_Energy_Bin_640 <= s_Energy_Bin_640 +'1';
		 Energy_Bin_Rdy_640 <= '1';
		else
		 s_Energy_Bin_640 <= s_Energy_Bin_640;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_640 <= '0';
      end if;
    end if;
  end process  Energy_Bin_640;    
  
  Energy_Bin_641 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_641   <=  (others =>'0');
		Energy_Bin_Rdy_641 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E641_C1_L and PEAK_C1 <= s_E641_C1_H and Bin_OR = '0') then
         s_Energy_Bin_641 <= s_Energy_Bin_641 +'1';
		 Energy_Bin_Rdy_641 <= '1';
		else
		 s_Energy_Bin_641 <= s_Energy_Bin_641;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_641 <= '0';
      end if;
    end if;
  end process  Energy_Bin_641;   
  
  Energy_Bin_642 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_642   <=  (others =>'0');
	    Energy_Bin_Rdy_642 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E642_C1_L and PEAK_C1 <= s_E642_C1_H and Bin_OR = '0') then
         s_Energy_Bin_642 <= s_Energy_Bin_642 +'1';
		 Energy_Bin_Rdy_642 <= '1';
		else
		 s_Energy_Bin_642 <= s_Energy_Bin_642;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_642 <= '0';
      end if;
    end if;
  end process  Energy_Bin_642;   
  
  Energy_Bin_643 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_643   <=  (others =>'0');
	    Energy_Bin_Rdy_643 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E643_C1_L and PEAK_C1 <= s_E643_C1_H and Bin_OR = '0') then
         s_Energy_Bin_643 <= s_Energy_Bin_643 +'1';
		 Energy_Bin_Rdy_643 <= '1';
		else
		 s_Energy_Bin_643 <= s_Energy_Bin_643;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_643 <= '0';
      end if;
    end if;
  end process  Energy_Bin_643;   
  
  Energy_Bin_644 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_644   <=  (others =>'0');
		Energy_Bin_Rdy_644 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E644_C1_L and PEAK_C1 <= s_E644_C1_H and Bin_OR = '0') then
         s_Energy_Bin_644 <= s_Energy_Bin_644 +'1';
		 Energy_Bin_Rdy_644 <= '1';
		else
		 s_Energy_Bin_644 <= s_Energy_Bin_644;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_644 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_644;   
 
 
  Energy_Bin_645 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_645   <=  (others =>'0');
		Energy_Bin_Rdy_645 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E645_C1_L and PEAK_C1 <= s_E645_C1_H and Bin_OR = '0') then
         s_Energy_Bin_645 <= s_Energy_Bin_645 +'1';
		 Energy_Bin_Rdy_645 <= '1';
		else
		 s_Energy_Bin_645 <= s_Energy_Bin_645;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_645 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_645;  
 
  
  Energy_Bin_646 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_646   <=  (others =>'0');
		Energy_Bin_Rdy_646 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E646_C1_L and PEAK_C1 <= s_E646_C1_H and Bin_OR = '0') then
         s_Energy_Bin_646 <= s_Energy_Bin_646 +'1';
		 Energy_Bin_Rdy_646 <= '1';
		else
		 s_Energy_Bin_646 <= s_Energy_Bin_646;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_646 <= '0';
      end if;
    end if;
  end process  Energy_Bin_646;   
  
 Energy_Bin_647 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_647   <=  (others =>'0');
		Energy_Bin_Rdy_647 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E647_C1_L and PEAK_C1 <= s_E647_C1_H and Bin_OR = '0') then
         s_Energy_Bin_647 <= s_Energy_Bin_647 +'1';
		 Energy_Bin_Rdy_647 <= '1';
		else
		 s_Energy_Bin_647 <= s_Energy_Bin_647;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_647 <= '0';
      end if;
    end if;
  end process  Energy_Bin_647;   
  
  Energy_Bin_648 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_648   <=  (others =>'0');
		Energy_Bin_Rdy_648 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E648_C1_L and PEAK_C1 <= s_E648_C1_H and Bin_OR = '0') then
         s_Energy_Bin_648 <= s_Energy_Bin_648 +'1';
		 Energy_Bin_Rdy_648 <= '1';
		else
		 s_Energy_Bin_648 <= s_Energy_Bin_648;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_648 <= '0';
      end if;
    end if;
  end process  Energy_Bin_648;   
  
  Energy_Bin_649 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_649   <=  (others =>'0');
		Energy_Bin_Rdy_649 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E649_C1_L and PEAK_C1 <= s_E649_C1_H and Bin_OR = '0') then
         s_Energy_Bin_649 <= s_Energy_Bin_649 +'1';
		 Energy_Bin_Rdy_649 <= '1';
		else
		 s_Energy_Bin_649 <= s_Energy_Bin_649;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_649 <= '0';
      end if;
    end if;
  end process  Energy_Bin_649;          
  
  
     Energy_Bin_650 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_650   <=  (others =>'0');
		Energy_Bin_Rdy_650 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E650_C1_L and PEAK_C1 <= s_E650_C1_H and Bin_OR = '0') then
         s_Energy_Bin_650 <= s_Energy_Bin_650 +'1';
		 Energy_Bin_Rdy_650 <= '1';
		else
		 s_Energy_Bin_650 <= s_Energy_Bin_650;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_650 <= '0';
      end if;
    end if;
  end process  Energy_Bin_650;    
  
  Energy_Bin_651 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_651   <=  (others =>'0');
		Energy_Bin_Rdy_651 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E651_C1_L and PEAK_C1 <= s_E651_C1_H and Bin_OR = '0') then
         s_Energy_Bin_651 <= s_Energy_Bin_651 +'1';
		 Energy_Bin_Rdy_651 <= '1';
		else
		 s_Energy_Bin_651 <= s_Energy_Bin_651;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_651 <= '0';
      end if;
    end if;
  end process  Energy_Bin_651;   
  
  Energy_Bin_652 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_652   <=  (others =>'0');
	    Energy_Bin_Rdy_652 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E652_C1_L and PEAK_C1 <= s_E652_C1_H and Bin_OR = '0') then
         s_Energy_Bin_652 <= s_Energy_Bin_652 +'1';
		 Energy_Bin_Rdy_652 <= '1';
		else
		 s_Energy_Bin_652 <= s_Energy_Bin_652;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_652 <= '0';
      end if;
    end if;
  end process  Energy_Bin_652;   
  
  Energy_Bin_653 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_653   <=  (others =>'0');
	    Energy_Bin_Rdy_653 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E653_C1_L and PEAK_C1 <= s_E653_C1_H and Bin_OR = '0') then
         s_Energy_Bin_653 <= s_Energy_Bin_653 +'1';
		 Energy_Bin_Rdy_653 <= '1';
		else
		 s_Energy_Bin_653 <= s_Energy_Bin_653;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_653 <= '0';
      end if;
    end if;
  end process  Energy_Bin_653;   
  
  Energy_Bin_654 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_654   <=  (others =>'0');
		Energy_Bin_Rdy_654 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E654_C1_L and PEAK_C1 <= s_E654_C1_H and Bin_OR = '0') then
         s_Energy_Bin_654 <= s_Energy_Bin_654 +'1';
		 Energy_Bin_Rdy_654 <= '1';
		else
		 s_Energy_Bin_654 <= s_Energy_Bin_654;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_654 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_654;   
 
 
  Energy_Bin_655 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_655   <=  (others =>'0');
		Energy_Bin_Rdy_655 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E655_C1_L and PEAK_C1 <= s_E655_C1_H and Bin_OR = '0') then
         s_Energy_Bin_655 <= s_Energy_Bin_655 +'1';
		 Energy_Bin_Rdy_655 <= '1';
		else
		 s_Energy_Bin_655 <= s_Energy_Bin_655;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_655 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_655;  
 
  
  Energy_Bin_656 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_656   <=  (others =>'0');
		Energy_Bin_Rdy_656 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E656_C1_L and PEAK_C1 <= s_E656_C1_H and Bin_OR = '0') then
         s_Energy_Bin_656 <= s_Energy_Bin_656 +'1';
		 Energy_Bin_Rdy_656 <= '1';
		else
		 s_Energy_Bin_656 <= s_Energy_Bin_656;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_656 <= '0';
      end if;
    end if;
  end process  Energy_Bin_656;   
  
 Energy_Bin_657 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_657   <=  (others =>'0');
		Energy_Bin_Rdy_657 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E657_C1_L and PEAK_C1 <= s_E657_C1_H and Bin_OR = '0') then
         s_Energy_Bin_657 <= s_Energy_Bin_657 +'1';
		 Energy_Bin_Rdy_657 <= '1';
		else
		 s_Energy_Bin_657 <= s_Energy_Bin_657;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_657 <= '0';
      end if;
    end if;
  end process  Energy_Bin_657;   
  
  Energy_Bin_658 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_658   <=  (others =>'0');
		Energy_Bin_Rdy_658 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E658_C1_L and PEAK_C1 <= s_E658_C1_H and Bin_OR = '0') then
         s_Energy_Bin_658 <= s_Energy_Bin_658 +'1';
		 Energy_Bin_Rdy_658 <= '1';
		else
		 s_Energy_Bin_658 <= s_Energy_Bin_658;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_658 <= '0';
      end if;
    end if;
  end process  Energy_Bin_658;   
  
  Energy_Bin_659 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_659   <=  (others =>'0');
		Energy_Bin_Rdy_659 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E659_C1_L and PEAK_C1 <= s_E659_C1_H and Bin_OR = '0') then
         s_Energy_Bin_659 <= s_Energy_Bin_659 +'1';
		 Energy_Bin_Rdy_659 <= '1';
		else
		 s_Energy_Bin_659 <= s_Energy_Bin_659;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_659 <= '0';
      end if;
    end if;
  end process  Energy_Bin_659;           
  
     Energy_Bin_660 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_660   <=  (others =>'0');
		Energy_Bin_Rdy_660 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E660_C1_L and PEAK_C1 <= s_E660_C1_H and Bin_OR = '0') then
         s_Energy_Bin_660 <= s_Energy_Bin_660 +'1';
		 Energy_Bin_Rdy_660 <= '1';
		else
		 s_Energy_Bin_660 <= s_Energy_Bin_660;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_660 <= '0';
      end if;
    end if;
  end process  Energy_Bin_660;    
  
  Energy_Bin_661 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_661   <=  (others =>'0');
		Energy_Bin_Rdy_661 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E661_C1_L and PEAK_C1 <= s_E661_C1_H and Bin_OR = '0') then
         s_Energy_Bin_661 <= s_Energy_Bin_661 +'1';
		 Energy_Bin_Rdy_661 <= '1';
		else
		 s_Energy_Bin_661 <= s_Energy_Bin_661;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_661 <= '0';
      end if;
    end if;
  end process  Energy_Bin_661;   
  
  Energy_Bin_662 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_662   <=  (others =>'0');
	    Energy_Bin_Rdy_662 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E662_C1_L and PEAK_C1 <= s_E662_C1_H and Bin_OR = '0') then
         s_Energy_Bin_662 <= s_Energy_Bin_662 +'1';
		 Energy_Bin_Rdy_662 <= '1';
		else
		 s_Energy_Bin_662 <= s_Energy_Bin_662;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_662 <= '0';
      end if;
    end if;
  end process  Energy_Bin_662;   
  
  Energy_Bin_663 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_663   <=  (others =>'0');
	    Energy_Bin_Rdy_663 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E663_C1_L and PEAK_C1 <= s_E663_C1_H and Bin_OR = '0') then
         s_Energy_Bin_663 <= s_Energy_Bin_663 +'1';
		 Energy_Bin_Rdy_663 <= '1';
		else
		 s_Energy_Bin_663 <= s_Energy_Bin_663;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_663 <= '0';
      end if;
    end if;
  end process  Energy_Bin_663;   
  
  Energy_Bin_664 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_664   <=  (others =>'0');
		Energy_Bin_Rdy_664 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E664_C1_L and PEAK_C1 <= s_E664_C1_H and Bin_OR = '0') then
         s_Energy_Bin_664 <= s_Energy_Bin_664 +'1';
		 Energy_Bin_Rdy_664 <= '1';
		else
		 s_Energy_Bin_664 <= s_Energy_Bin_664;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_664 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_664;   
 
 
  Energy_Bin_665 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_665   <=  (others =>'0');
		Energy_Bin_Rdy_665 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E665_C1_L and PEAK_C1 <= s_E665_C1_H and Bin_OR = '0') then
         s_Energy_Bin_665 <= s_Energy_Bin_665 +'1';
		 Energy_Bin_Rdy_665 <= '1';
		else
		 s_Energy_Bin_665 <= s_Energy_Bin_665;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_665 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_665;  
 
  
  Energy_Bin_666 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_666   <=  (others =>'0');
		Energy_Bin_Rdy_666 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E666_C1_L and PEAK_C1 <= s_E666_C1_H and Bin_OR = '0') then
         s_Energy_Bin_666 <= s_Energy_Bin_666 +'1';
		 Energy_Bin_Rdy_666 <= '1';
		else
		 s_Energy_Bin_666 <= s_Energy_Bin_666;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_666 <= '0';
      end if;
    end if;
  end process  Energy_Bin_666;   
  
 Energy_Bin_667 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_667   <=  (others =>'0');
		Energy_Bin_Rdy_667 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E667_C1_L and PEAK_C1 <= s_E667_C1_H and Bin_OR = '0') then
         s_Energy_Bin_667 <= s_Energy_Bin_667 +'1';
		 Energy_Bin_Rdy_667 <= '1';
		else
		 s_Energy_Bin_667 <= s_Energy_Bin_667;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_667 <= '0';
      end if;
    end if;
  end process  Energy_Bin_667;   
  
  Energy_Bin_668 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_668   <=  (others =>'0');
		Energy_Bin_Rdy_668 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E668_C1_L and PEAK_C1 <= s_E668_C1_H and Bin_OR = '0') then
         s_Energy_Bin_668 <= s_Energy_Bin_668 +'1';
		 Energy_Bin_Rdy_668 <= '1';
		else
		 s_Energy_Bin_668 <= s_Energy_Bin_668;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_668 <= '0';
      end if;
    end if;
  end process  Energy_Bin_668;   
  
  Energy_Bin_669 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_669   <=  (others =>'0');
		Energy_Bin_Rdy_669 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E669_C1_L and PEAK_C1 <= s_E669_C1_H and Bin_OR = '0') then
         s_Energy_Bin_669 <= s_Energy_Bin_669 +'1';
		 Energy_Bin_Rdy_669 <= '1';
		else
		 s_Energy_Bin_669 <= s_Energy_Bin_669;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_669 <= '0';
      end if;
    end if;
  end process  Energy_Bin_669;         
  
     Energy_Bin_670 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_670   <=  (others =>'0');
		Energy_Bin_Rdy_670 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E670_C1_L and PEAK_C1 <= s_E670_C1_H and Bin_OR = '0') then
         s_Energy_Bin_670 <= s_Energy_Bin_670 +'1';
		 Energy_Bin_Rdy_670 <= '1';
		else
		 s_Energy_Bin_670 <= s_Energy_Bin_670;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_670 <= '0';
      end if;
    end if;
  end process  Energy_Bin_670;    
  
  Energy_Bin_671 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_671   <=  (others =>'0');
		Energy_Bin_Rdy_671 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E671_C1_L and PEAK_C1 <= s_E671_C1_H and Bin_OR = '0') then
         s_Energy_Bin_671 <= s_Energy_Bin_671 +'1';
		 Energy_Bin_Rdy_671 <= '1';
		else
		 s_Energy_Bin_671 <= s_Energy_Bin_671;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_671 <= '0';
      end if;
    end if;
  end process  Energy_Bin_671;   
  
  Energy_Bin_672 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_672   <=  (others =>'0');
	    Energy_Bin_Rdy_672 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E672_C1_L and PEAK_C1 <= s_E672_C1_H and Bin_OR = '0') then
         s_Energy_Bin_672 <= s_Energy_Bin_672 +'1';
		 Energy_Bin_Rdy_672 <= '1';
		else
		 s_Energy_Bin_672 <= s_Energy_Bin_672;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_672 <= '0';
      end if;
    end if;
  end process  Energy_Bin_672;   
  
  Energy_Bin_673 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_673   <=  (others =>'0');
	    Energy_Bin_Rdy_673 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E673_C1_L and PEAK_C1 <= s_E673_C1_H and Bin_OR = '0') then
         s_Energy_Bin_673 <= s_Energy_Bin_673 +'1';
		 Energy_Bin_Rdy_673 <= '1';
		else
		 s_Energy_Bin_673 <= s_Energy_Bin_673;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_673 <= '0';
      end if;
    end if;
  end process  Energy_Bin_673;   
  
  Energy_Bin_674 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_674   <=  (others =>'0');
		Energy_Bin_Rdy_674 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E674_C1_L and PEAK_C1 <= s_E674_C1_H and Bin_OR = '0') then
         s_Energy_Bin_674 <= s_Energy_Bin_674 +'1';
		 Energy_Bin_Rdy_674 <= '1';
		else
		 s_Energy_Bin_674 <= s_Energy_Bin_674;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_674 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_674;   
 
 
  Energy_Bin_675 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_675   <=  (others =>'0');
		Energy_Bin_Rdy_675 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E675_C1_L and PEAK_C1 <= s_E675_C1_H and Bin_OR = '0') then
         s_Energy_Bin_675 <= s_Energy_Bin_675 +'1';
		 Energy_Bin_Rdy_675 <= '1';
		else
		 s_Energy_Bin_675 <= s_Energy_Bin_675;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_675 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_675;  
 
  
  Energy_Bin_676 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_676   <=  (others =>'0');
		Energy_Bin_Rdy_676 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E676_C1_L and PEAK_C1 <= s_E676_C1_H and Bin_OR = '0') then
         s_Energy_Bin_676 <= s_Energy_Bin_676 +'1';
		 Energy_Bin_Rdy_676 <= '1';
		else
		 s_Energy_Bin_676 <= s_Energy_Bin_676;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_676 <= '0';
      end if;
    end if;
  end process  Energy_Bin_676;   
  
 Energy_Bin_677 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_677   <=  (others =>'0');
		Energy_Bin_Rdy_677 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E677_C1_L and PEAK_C1 <= s_E677_C1_H and Bin_OR = '0') then
         s_Energy_Bin_677 <= s_Energy_Bin_677 +'1';
		 Energy_Bin_Rdy_677 <= '1';
		else
		 s_Energy_Bin_677 <= s_Energy_Bin_677;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_677 <= '0';
      end if;
    end if;
  end process  Energy_Bin_677;   
  
  Energy_Bin_678 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_678   <=  (others =>'0');
		Energy_Bin_Rdy_678 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E678_C1_L and PEAK_C1 <= s_E678_C1_H and Bin_OR = '0') then
         s_Energy_Bin_678 <= s_Energy_Bin_678 +'1';
		 Energy_Bin_Rdy_678 <= '1';
		else
		 s_Energy_Bin_678 <= s_Energy_Bin_678;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_678 <= '0';
      end if;
    end if;
  end process  Energy_Bin_678;   
  
  Energy_Bin_679 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_679   <=  (others =>'0');
		Energy_Bin_Rdy_679 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E679_C1_L and PEAK_C1 <= s_E679_C1_H and Bin_OR = '0') then
         s_Energy_Bin_679 <= s_Energy_Bin_679 +'1';
		 Energy_Bin_Rdy_679 <= '1';
		else
		 s_Energy_Bin_679 <= s_Energy_Bin_679;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_679 <= '0';
      end if;
    end if;
  end process  Energy_Bin_679;       
  
     Energy_Bin_680 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_680   <=  (others =>'0');
		Energy_Bin_Rdy_680 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E680_C1_L and PEAK_C1 <= s_E680_C1_H and Bin_OR = '0') then
         s_Energy_Bin_680 <= s_Energy_Bin_680 +'1';
		 Energy_Bin_Rdy_680 <= '1';
		else
		 s_Energy_Bin_680 <= s_Energy_Bin_680;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_680 <= '0';
      end if;
    end if;
  end process  Energy_Bin_680;    
  
  Energy_Bin_681 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_681   <=  (others =>'0');
		Energy_Bin_Rdy_681 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E681_C1_L and PEAK_C1 <= s_E681_C1_H and Bin_OR = '0') then
         s_Energy_Bin_681 <= s_Energy_Bin_681 +'1';
		 Energy_Bin_Rdy_681 <= '1';
		else
		 s_Energy_Bin_681 <= s_Energy_Bin_681;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_681 <= '0';
      end if;
    end if;
  end process  Energy_Bin_681;   
  
  Energy_Bin_682 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_682   <=  (others =>'0');
	    Energy_Bin_Rdy_682 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E682_C1_L and PEAK_C1 <= s_E682_C1_H and Bin_OR = '0') then
         s_Energy_Bin_682 <= s_Energy_Bin_682 +'1';
		 Energy_Bin_Rdy_682 <= '1';
		else
		 s_Energy_Bin_682 <= s_Energy_Bin_682;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_682 <= '0';
      end if;
    end if;
  end process  Energy_Bin_682;   
  
  Energy_Bin_683 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_683   <=  (others =>'0');
	    Energy_Bin_Rdy_683 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E683_C1_L and PEAK_C1 <= s_E683_C1_H and Bin_OR = '0') then
         s_Energy_Bin_683 <= s_Energy_Bin_683 +'1';
		 Energy_Bin_Rdy_683 <= '1';
		else
		 s_Energy_Bin_683 <= s_Energy_Bin_683;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_683 <= '0';
      end if;
    end if;
  end process  Energy_Bin_683;   
  
  Energy_Bin_684 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_684   <=  (others =>'0');
		Energy_Bin_Rdy_684 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E684_C1_L and PEAK_C1 <= s_E684_C1_H and Bin_OR = '0') then
         s_Energy_Bin_684 <= s_Energy_Bin_684 +'1';
		 Energy_Bin_Rdy_684 <= '1';
		else
		 s_Energy_Bin_684 <= s_Energy_Bin_684;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_684 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_684;   
 
 
  Energy_Bin_685 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_685   <=  (others =>'0');
		Energy_Bin_Rdy_685 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E685_C1_L and PEAK_C1 <= s_E685_C1_H and Bin_OR = '0') then
         s_Energy_Bin_685 <= s_Energy_Bin_685 +'1';
		 Energy_Bin_Rdy_685 <= '1';
		else
		 s_Energy_Bin_685 <= s_Energy_Bin_685;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_685 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_685;  
 
  
  Energy_Bin_686 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_686   <=  (others =>'0');
		Energy_Bin_Rdy_686 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E686_C1_L and PEAK_C1 <= s_E686_C1_H and Bin_OR = '0') then
         s_Energy_Bin_686 <= s_Energy_Bin_686 +'1';
		 Energy_Bin_Rdy_686 <= '1';
		else
		 s_Energy_Bin_686 <= s_Energy_Bin_686;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_686 <= '0';
      end if;
    end if;
  end process  Energy_Bin_686;   
  
 Energy_Bin_687 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_687   <=  (others =>'0');
		Energy_Bin_Rdy_687 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E687_C1_L and PEAK_C1 <= s_E687_C1_H and Bin_OR = '0') then
         s_Energy_Bin_687 <= s_Energy_Bin_687 +'1';
		 Energy_Bin_Rdy_687 <= '1';
		else
		 s_Energy_Bin_687 <= s_Energy_Bin_687;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_687 <= '0';
      end if;
    end if;
  end process  Energy_Bin_687;   
  
  Energy_Bin_688 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_688   <=  (others =>'0');
		Energy_Bin_Rdy_688 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E688_C1_L and PEAK_C1 <= s_E688_C1_H and Bin_OR = '0') then
         s_Energy_Bin_688 <= s_Energy_Bin_688 +'1';
		 Energy_Bin_Rdy_688 <= '1';
		else
		 s_Energy_Bin_688 <= s_Energy_Bin_688;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_688 <= '0';
      end if;
    end if;
  end process  Energy_Bin_688;   
  
  Energy_Bin_689 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_689   <=  (others =>'0');
		Energy_Bin_Rdy_689 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E689_C1_L and PEAK_C1 <= s_E689_C1_H and Bin_OR = '0') then
         s_Energy_Bin_689 <= s_Energy_Bin_689 +'1';
		 Energy_Bin_Rdy_689 <= '1';
		else
		 s_Energy_Bin_689 <= s_Energy_Bin_689;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_689 <= '0';
      end if;
    end if;
  end process  Energy_Bin_689;      
  
     Energy_Bin_690 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_690   <=  (others =>'0');
		Energy_Bin_Rdy_690 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E690_C1_L and PEAK_C1 <= s_E690_C1_H and Bin_OR = '0') then
         s_Energy_Bin_690 <= s_Energy_Bin_690 +'1';
		 Energy_Bin_Rdy_690 <= '1';
		else
		 s_Energy_Bin_690 <= s_Energy_Bin_690;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_690 <= '0';
      end if;
    end if;
  end process  Energy_Bin_690;    
  
  Energy_Bin_691 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_691   <=  (others =>'0');
		Energy_Bin_Rdy_691 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E691_C1_L and PEAK_C1 <= s_E691_C1_H and Bin_OR = '0') then
         s_Energy_Bin_691 <= s_Energy_Bin_691 +'1';
		 Energy_Bin_Rdy_691 <= '1';
		else
		 s_Energy_Bin_691 <= s_Energy_Bin_691;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_691 <= '0';
      end if;
    end if;
  end process  Energy_Bin_691;   
  
  Energy_Bin_692 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_692   <=  (others =>'0');
	    Energy_Bin_Rdy_692 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E692_C1_L and PEAK_C1 <= s_E692_C1_H and Bin_OR = '0') then
         s_Energy_Bin_692 <= s_Energy_Bin_692 +'1';
		 Energy_Bin_Rdy_692 <= '1';
		else
		 s_Energy_Bin_692 <= s_Energy_Bin_692;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_692 <= '0';
      end if;
    end if;
  end process  Energy_Bin_692;   
  
  Energy_Bin_693 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_693   <=  (others =>'0');
	    Energy_Bin_Rdy_693 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E693_C1_L and PEAK_C1 <= s_E693_C1_H and Bin_OR = '0') then
         s_Energy_Bin_693 <= s_Energy_Bin_693 +'1';
		 Energy_Bin_Rdy_693 <= '1';
		else
		 s_Energy_Bin_693 <= s_Energy_Bin_693;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_693 <= '0';
      end if;
    end if;
  end process  Energy_Bin_693;   
  
  Energy_Bin_694 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_694   <=  (others =>'0');
		Energy_Bin_Rdy_694 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E694_C1_L and PEAK_C1 <= s_E694_C1_H and Bin_OR = '0') then
         s_Energy_Bin_694 <= s_Energy_Bin_694 +'1';
		 Energy_Bin_Rdy_694 <= '1';
		else
		 s_Energy_Bin_694 <= s_Energy_Bin_694;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_694 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_694;   
 
 
  Energy_Bin_695 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_695   <=  (others =>'0');
		Energy_Bin_Rdy_695 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E695_C1_L and PEAK_C1 <= s_E695_C1_H and Bin_OR = '0') then
         s_Energy_Bin_695 <= s_Energy_Bin_695 +'1';
		 Energy_Bin_Rdy_695 <= '1';
		else
		 s_Energy_Bin_695 <= s_Energy_Bin_695;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_695 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_695;  
 
  
  Energy_Bin_696 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_696   <=  (others =>'0');
		Energy_Bin_Rdy_696 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E696_C1_L and PEAK_C1 <= s_E696_C1_H and Bin_OR = '0') then
         s_Energy_Bin_696 <= s_Energy_Bin_696 +'1';
		 Energy_Bin_Rdy_696 <= '1';
		else
		 s_Energy_Bin_696 <= s_Energy_Bin_696;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_696 <= '0';
      end if;
    end if;
  end process  Energy_Bin_696;   
  
 Energy_Bin_697 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_697   <=  (others =>'0');
		Energy_Bin_Rdy_697 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E697_C1_L and PEAK_C1 <= s_E697_C1_H and Bin_OR = '0') then
         s_Energy_Bin_697 <= s_Energy_Bin_697 +'1';
		 Energy_Bin_Rdy_697 <= '1';
		else
		 s_Energy_Bin_697 <= s_Energy_Bin_697;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_697 <= '0';
      end if;
    end if;
  end process  Energy_Bin_697;   
  
  Energy_Bin_698 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_698   <=  (others =>'0');
		Energy_Bin_Rdy_698 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E698_C1_L and PEAK_C1 <= s_E698_C1_H and Bin_OR = '0') then
         s_Energy_Bin_698 <= s_Energy_Bin_698 +'1';
		 Energy_Bin_Rdy_698 <= '1';
		else
		 s_Energy_Bin_698 <= s_Energy_Bin_698;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_698 <= '0';
      end if;
    end if;
  end process  Energy_Bin_698;   
  
  Energy_Bin_699 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_699   <=  (others =>'0');
		Energy_Bin_Rdy_699 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E699_C1_L and PEAK_C1 <= s_E699_C1_H and Bin_OR = '0') then
         s_Energy_Bin_699 <= s_Energy_Bin_699 +'1';
		 Energy_Bin_Rdy_699 <= '1';
		else
		 s_Energy_Bin_699 <= s_Energy_Bin_699;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_699 <= '0';
      end if;
    end if;
  end process  Energy_Bin_699;   

    Energy_Bin_700 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_700   <=  (others =>'0');
		Energy_Bin_Rdy_700 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E700_C1_L and PEAK_C1 <= s_E700_C1_H and Bin_OR = '0') then
         s_Energy_Bin_700 <= s_Energy_Bin_700 +'1';
		 Energy_Bin_Rdy_700 <= '1';
		else
		 s_Energy_Bin_700 <= s_Energy_Bin_700;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_700 <= '0';
      end if;
    end if;
  end process  Energy_Bin_700;    
  
  Energy_Bin_701 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_701   <=  (others =>'0');
		Energy_Bin_Rdy_701 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E701_C1_L and PEAK_C1 <= s_E701_C1_H and Bin_OR = '0') then
         s_Energy_Bin_701 <= s_Energy_Bin_701 +'1';
		 Energy_Bin_Rdy_701 <= '1';
		else
		 s_Energy_Bin_701 <= s_Energy_Bin_701;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_701 <= '0';
      end if;
    end if;
  end process  Energy_Bin_701;   
  
  Energy_Bin_702 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_702   <=  (others =>'0');
	    Energy_Bin_Rdy_702 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E702_C1_L and PEAK_C1 <= s_E702_C1_H and Bin_OR = '0') then
         s_Energy_Bin_702 <= s_Energy_Bin_702 +'1';
		 Energy_Bin_Rdy_702 <= '1';
		else
		 s_Energy_Bin_702 <= s_Energy_Bin_702;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_702 <= '0';
      end if;
    end if;
  end process  Energy_Bin_702;   
  
  Energy_Bin_703 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_703   <=  (others =>'0');
	    Energy_Bin_Rdy_703 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E703_C1_L and PEAK_C1 <= s_E703_C1_H and Bin_OR = '0') then
         s_Energy_Bin_703 <= s_Energy_Bin_703 +'1';
		 Energy_Bin_Rdy_703 <= '1';
		else
		 s_Energy_Bin_703 <= s_Energy_Bin_703;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_703 <= '0';
      end if;
    end if;
  end process  Energy_Bin_703;   
  
  Energy_Bin_704 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_704   <=  (others =>'0');
		Energy_Bin_Rdy_704 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E704_C1_L and PEAK_C1 <= s_E704_C1_H and Bin_OR = '0') then
         s_Energy_Bin_704 <= s_Energy_Bin_704 +'1';
		 Energy_Bin_Rdy_704 <= '1';
		else
		 s_Energy_Bin_704 <= s_Energy_Bin_704;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_704 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_704;   
 
 
  Energy_Bin_705 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_705   <=  (others =>'0');
		Energy_Bin_Rdy_705 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E705_C1_L and PEAK_C1 <= s_E705_C1_H and Bin_OR = '0') then
         s_Energy_Bin_705 <= s_Energy_Bin_705 +'1';
		 Energy_Bin_Rdy_705 <= '1';
		else
		 s_Energy_Bin_705 <= s_Energy_Bin_705;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_705 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_705;  
 
  
  Energy_Bin_706 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_706   <=  (others =>'0');
		Energy_Bin_Rdy_706 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E706_C1_L and PEAK_C1 <= s_E706_C1_H and Bin_OR = '0') then
         s_Energy_Bin_706 <= s_Energy_Bin_706 +'1';
		 Energy_Bin_Rdy_706 <= '1';
		else
		 s_Energy_Bin_706 <= s_Energy_Bin_706;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_706 <= '0';
      end if;
    end if;
  end process  Energy_Bin_706;   
  
 Energy_Bin_707 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_707   <=  (others =>'0');
		Energy_Bin_Rdy_707 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E707_C1_L and PEAK_C1 <= s_E707_C1_H and Bin_OR = '0') then
         s_Energy_Bin_707 <= s_Energy_Bin_707 +'1';
		 Energy_Bin_Rdy_707 <= '1';
		else
		 s_Energy_Bin_707 <= s_Energy_Bin_707;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_707 <= '0';
      end if;
    end if;
  end process  Energy_Bin_707;   
  
  Energy_Bin_708 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_708   <=  (others =>'0');
		Energy_Bin_Rdy_708 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E708_C1_L and PEAK_C1 <= s_E708_C1_H and Bin_OR = '0') then
         s_Energy_Bin_708 <= s_Energy_Bin_708 +'1';
		 Energy_Bin_Rdy_708 <= '1';
		else
		 s_Energy_Bin_708 <= s_Energy_Bin_708;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_708 <= '0';
      end if;
    end if;
  end process  Energy_Bin_708;   
  
  Energy_Bin_709 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_709   <=  (others =>'0');
		Energy_Bin_Rdy_709 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E709_C1_L and PEAK_C1 <= s_E709_C1_H and Bin_OR = '0') then
         s_Energy_Bin_709 <= s_Energy_Bin_709 +'1';
		 Energy_Bin_Rdy_709 <= '1';
		else
		 s_Energy_Bin_709 <= s_Energy_Bin_709;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_709 <= '0';
      end if;
    end if;
  end process  Energy_Bin_709;      
  
     Energy_Bin_710 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_710   <=  (others =>'0');
		Energy_Bin_Rdy_710 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E710_C1_L and PEAK_C1 <= s_E710_C1_H and Bin_OR = '0') then
         s_Energy_Bin_710 <= s_Energy_Bin_710 +'1';
		 Energy_Bin_Rdy_710 <= '1';
		else
		 s_Energy_Bin_710 <= s_Energy_Bin_710;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_710 <= '0';
      end if;
    end if;
  end process  Energy_Bin_710;    
  
  Energy_Bin_711 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_711   <=  (others =>'0');
		Energy_Bin_Rdy_711 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E711_C1_L and PEAK_C1 <= s_E711_C1_H and Bin_OR = '0') then
         s_Energy_Bin_711 <= s_Energy_Bin_711 +'1';
		 Energy_Bin_Rdy_711 <= '1';
		else
		 s_Energy_Bin_711 <= s_Energy_Bin_711;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_711 <= '0';
      end if;
    end if;
  end process  Energy_Bin_711;   
  
  Energy_Bin_712 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_712   <=  (others =>'0');
	    Energy_Bin_Rdy_712 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E712_C1_L and PEAK_C1 <= s_E712_C1_H and Bin_OR = '0') then
         s_Energy_Bin_712 <= s_Energy_Bin_712 +'1';
		 Energy_Bin_Rdy_712 <= '1';
		else
		 s_Energy_Bin_712 <= s_Energy_Bin_712;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_712 <= '0';
      end if;
    end if;
  end process  Energy_Bin_712;   
  
  Energy_Bin_713 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_713   <=  (others =>'0');
	    Energy_Bin_Rdy_713 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E713_C1_L and PEAK_C1 <= s_E713_C1_H and Bin_OR = '0') then
         s_Energy_Bin_713 <= s_Energy_Bin_713 +'1';
		 Energy_Bin_Rdy_713 <= '1';
		else
		 s_Energy_Bin_713 <= s_Energy_Bin_713;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_713 <= '0';
      end if;
    end if;
  end process  Energy_Bin_713;   
  
  Energy_Bin_714 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_714   <=  (others =>'0');
		Energy_Bin_Rdy_714 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E714_C1_L and PEAK_C1 <= s_E714_C1_H and Bin_OR = '0') then
         s_Energy_Bin_714 <= s_Energy_Bin_714 +'1';
		 Energy_Bin_Rdy_714 <= '1';
		else
		 s_Energy_Bin_714 <= s_Energy_Bin_714;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_714 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_714;   
 
 
  Energy_Bin_715 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_715   <=  (others =>'0');
		Energy_Bin_Rdy_715 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E715_C1_L and PEAK_C1 <= s_E715_C1_H and Bin_OR = '0') then
         s_Energy_Bin_715 <= s_Energy_Bin_715 +'1';
		 Energy_Bin_Rdy_715 <= '1';
		else
		 s_Energy_Bin_715 <= s_Energy_Bin_715;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_715 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_715;  
 
  
  Energy_Bin_716 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_716   <=  (others =>'0');
		Energy_Bin_Rdy_716 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E716_C1_L and PEAK_C1 <= s_E716_C1_H and Bin_OR = '0') then
         s_Energy_Bin_716 <= s_Energy_Bin_716 +'1';
		 Energy_Bin_Rdy_716 <= '1';
		else
		 s_Energy_Bin_716 <= s_Energy_Bin_716;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_716 <= '0';
      end if;
    end if;
  end process  Energy_Bin_716;   
  
 Energy_Bin_717 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_717   <=  (others =>'0');
		Energy_Bin_Rdy_717 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E717_C1_L and PEAK_C1 <= s_E717_C1_H and Bin_OR = '0') then
         s_Energy_Bin_717 <= s_Energy_Bin_717 +'1';
		 Energy_Bin_Rdy_717 <= '1';
		else
		 s_Energy_Bin_717 <= s_Energy_Bin_717;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_717 <= '0';
      end if;
    end if;
  end process  Energy_Bin_717;   
  
  Energy_Bin_718 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_718   <=  (others =>'0');
		Energy_Bin_Rdy_718 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E718_C1_L and PEAK_C1 <= s_E718_C1_H and Bin_OR = '0') then
         s_Energy_Bin_718 <= s_Energy_Bin_718 +'1';
		 Energy_Bin_Rdy_718 <= '1';
		else
		 s_Energy_Bin_718 <= s_Energy_Bin_718;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_718 <= '0';
      end if;
    end if;
  end process  Energy_Bin_718;   
  
  Energy_Bin_719 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_719   <=  (others =>'0');
		Energy_Bin_Rdy_719 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E719_C1_L and PEAK_C1 <= s_E719_C1_H and Bin_OR = '0') then
         s_Energy_Bin_719 <= s_Energy_Bin_719 +'1';
		 Energy_Bin_Rdy_719 <= '1';
		else
		 s_Energy_Bin_719 <= s_Energy_Bin_719;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_719 <= '0';
      end if;
    end if;
  end process  Energy_Bin_719;       
  
     Energy_Bin_720 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_720   <=  (others =>'0');
		Energy_Bin_Rdy_720 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E720_C1_L and PEAK_C1 <= s_E720_C1_H and Bin_OR = '0') then
         s_Energy_Bin_720 <= s_Energy_Bin_720 +'1';
		 Energy_Bin_Rdy_720 <= '1';
		else
		 s_Energy_Bin_720 <= s_Energy_Bin_720;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_720 <= '0';
      end if;
    end if;
  end process  Energy_Bin_720;    
  
  Energy_Bin_721 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_721   <=  (others =>'0');
		Energy_Bin_Rdy_721 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E721_C1_L and PEAK_C1 <= s_E721_C1_H and Bin_OR = '0') then
         s_Energy_Bin_721 <= s_Energy_Bin_721 +'1';
		 Energy_Bin_Rdy_721 <= '1';
		else
		 s_Energy_Bin_721 <= s_Energy_Bin_721;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_721 <= '0';
      end if;
    end if;
  end process  Energy_Bin_721;   
  
  Energy_Bin_722 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_722   <=  (others =>'0');
	    Energy_Bin_Rdy_722 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E722_C1_L and PEAK_C1 <= s_E722_C1_H and Bin_OR = '0') then
         s_Energy_Bin_722 <= s_Energy_Bin_722 +'1';
		 Energy_Bin_Rdy_722 <= '1';
		else
		 s_Energy_Bin_722 <= s_Energy_Bin_722;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_722 <= '0';
      end if;
    end if;
  end process  Energy_Bin_722;   
  
  Energy_Bin_723 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_723   <=  (others =>'0');
	    Energy_Bin_Rdy_723 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E723_C1_L and PEAK_C1 <= s_E723_C1_H and Bin_OR = '0') then
         s_Energy_Bin_723 <= s_Energy_Bin_723 +'1';
		 Energy_Bin_Rdy_723 <= '1';
		else
		 s_Energy_Bin_723 <= s_Energy_Bin_723;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_723 <= '0';
      end if;
    end if;
  end process  Energy_Bin_723;   
  
  Energy_Bin_724 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_724   <=  (others =>'0');
		Energy_Bin_Rdy_724 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E724_C1_L and PEAK_C1 <= s_E724_C1_H and Bin_OR = '0') then
         s_Energy_Bin_724 <= s_Energy_Bin_724 +'1';
		 Energy_Bin_Rdy_724 <= '1';
		else
		 s_Energy_Bin_724 <= s_Energy_Bin_724;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_724 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_724;   
 
 
  Energy_Bin_725 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_725   <=  (others =>'0');
		Energy_Bin_Rdy_725 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E725_C1_L and PEAK_C1 <= s_E725_C1_H and Bin_OR = '0') then
         s_Energy_Bin_725 <= s_Energy_Bin_725 +'1';
		 Energy_Bin_Rdy_725 <= '1';
		else
		 s_Energy_Bin_725 <= s_Energy_Bin_725;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_725 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_725;  
 
  
  Energy_Bin_726 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_726   <=  (others =>'0');
		Energy_Bin_Rdy_726 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E726_C1_L and PEAK_C1 <= s_E726_C1_H and Bin_OR = '0') then
         s_Energy_Bin_726 <= s_Energy_Bin_726 +'1';
		 Energy_Bin_Rdy_726 <= '1';
		else
		 s_Energy_Bin_726 <= s_Energy_Bin_726;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_726 <= '0';
      end if;
    end if;
  end process  Energy_Bin_726;   
  
 Energy_Bin_727 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_727   <=  (others =>'0');
		Energy_Bin_Rdy_727 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E727_C1_L and PEAK_C1 <= s_E727_C1_H and Bin_OR = '0') then
         s_Energy_Bin_727 <= s_Energy_Bin_727 +'1';
		 Energy_Bin_Rdy_727 <= '1';
		else
		 s_Energy_Bin_727 <= s_Energy_Bin_727;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_727 <= '0';
      end if;
    end if;
  end process  Energy_Bin_727;   
  
  Energy_Bin_728 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_728   <=  (others =>'0');
		Energy_Bin_Rdy_728 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E728_C1_L and PEAK_C1 <= s_E728_C1_H and Bin_OR = '0') then
         s_Energy_Bin_728 <= s_Energy_Bin_728 +'1';
		 Energy_Bin_Rdy_728 <= '1';
		else
		 s_Energy_Bin_728 <= s_Energy_Bin_728;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_728 <= '0';
      end if;
    end if;
  end process  Energy_Bin_728;   
  
  Energy_Bin_729 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_729   <=  (others =>'0');
		Energy_Bin_Rdy_729 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E729_C1_L and PEAK_C1 <= s_E729_C1_H and Bin_OR = '0') then
         s_Energy_Bin_729 <= s_Energy_Bin_729 +'1';
		 Energy_Bin_Rdy_729 <= '1';
		else
		 s_Energy_Bin_729 <= s_Energy_Bin_729;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_729 <= '0';
      end if;
    end if;
  end process  Energy_Bin_729;        
  
     Energy_Bin_730 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_730   <=  (others =>'0');
		Energy_Bin_Rdy_730 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E730_C1_L and PEAK_C1 <= s_E730_C1_H and Bin_OR = '0') then
         s_Energy_Bin_730 <= s_Energy_Bin_730 +'1';
		 Energy_Bin_Rdy_730 <= '1';
		else
		 s_Energy_Bin_730 <= s_Energy_Bin_730;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_730 <= '0';
      end if;
    end if;
  end process  Energy_Bin_730;    
  
  Energy_Bin_731 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_731   <=  (others =>'0');
		Energy_Bin_Rdy_731 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E731_C1_L and PEAK_C1 <= s_E731_C1_H and Bin_OR = '0') then
         s_Energy_Bin_731 <= s_Energy_Bin_731 +'1';
		 Energy_Bin_Rdy_731 <= '1';
		else
		 s_Energy_Bin_731 <= s_Energy_Bin_731;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_731 <= '0';
      end if;
    end if;
  end process  Energy_Bin_731;   
  
  Energy_Bin_732 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_732   <=  (others =>'0');
	    Energy_Bin_Rdy_732 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E732_C1_L and PEAK_C1 <= s_E732_C1_H and Bin_OR = '0') then
         s_Energy_Bin_732 <= s_Energy_Bin_732 +'1';
		 Energy_Bin_Rdy_732 <= '1';
		else
		 s_Energy_Bin_732 <= s_Energy_Bin_732;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_732 <= '0';
      end if;
    end if;
  end process  Energy_Bin_732;   
  
  Energy_Bin_733 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_733   <=  (others =>'0');
	    Energy_Bin_Rdy_733 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E733_C1_L and PEAK_C1 <= s_E733_C1_H and Bin_OR = '0') then
         s_Energy_Bin_733 <= s_Energy_Bin_733 +'1';
		 Energy_Bin_Rdy_733 <= '1';
		else
		 s_Energy_Bin_733 <= s_Energy_Bin_733;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_733 <= '0';
      end if;
    end if;
  end process  Energy_Bin_733;   
  
  Energy_Bin_734 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_734   <=  (others =>'0');
		Energy_Bin_Rdy_734 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E734_C1_L and PEAK_C1 <= s_E734_C1_H and Bin_OR = '0') then
         s_Energy_Bin_734 <= s_Energy_Bin_734 +'1';
		 Energy_Bin_Rdy_734 <= '1';
		else
		 s_Energy_Bin_734 <= s_Energy_Bin_734;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_734 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_734;   
 
 
  Energy_Bin_735 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_735   <=  (others =>'0');
		Energy_Bin_Rdy_735 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E735_C1_L and PEAK_C1 <= s_E735_C1_H and Bin_OR = '0') then
         s_Energy_Bin_735 <= s_Energy_Bin_735 +'1';
		 Energy_Bin_Rdy_735 <= '1';
		else
		 s_Energy_Bin_735 <= s_Energy_Bin_735;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_735 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_735;  
 
  
  Energy_Bin_736 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_736   <=  (others =>'0');
		Energy_Bin_Rdy_736 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E736_C1_L and PEAK_C1 <= s_E736_C1_H and Bin_OR = '0') then
         s_Energy_Bin_736 <= s_Energy_Bin_736 +'1';
		 Energy_Bin_Rdy_736 <= '1';
		else
		 s_Energy_Bin_736 <= s_Energy_Bin_736;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_736 <= '0';
      end if;
    end if;
  end process  Energy_Bin_736;   
  
 Energy_Bin_737 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_737   <=  (others =>'0');
		Energy_Bin_Rdy_737 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E737_C1_L and PEAK_C1 <= s_E737_C1_H and Bin_OR = '0') then
         s_Energy_Bin_737 <= s_Energy_Bin_737 +'1';
		 Energy_Bin_Rdy_737 <= '1';
		else
		 s_Energy_Bin_737 <= s_Energy_Bin_737;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_737 <= '0';
      end if;
    end if;
  end process  Energy_Bin_737;   
  
  Energy_Bin_738 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_738   <=  (others =>'0');
		Energy_Bin_Rdy_738 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E738_C1_L and PEAK_C1 <= s_E738_C1_H and Bin_OR = '0') then
         s_Energy_Bin_738 <= s_Energy_Bin_738 +'1';
		 Energy_Bin_Rdy_738 <= '1';
		else
		 s_Energy_Bin_738 <= s_Energy_Bin_738;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_738 <= '0';
      end if;
    end if;
  end process  Energy_Bin_738;   
  
  Energy_Bin_739 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_739   <=  (others =>'0');
		Energy_Bin_Rdy_739 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E739_C1_L and PEAK_C1 <= s_E739_C1_H and Bin_OR = '0') then
         s_Energy_Bin_739 <= s_Energy_Bin_739 +'1';
		 Energy_Bin_Rdy_739 <= '1';
		else
		 s_Energy_Bin_739 <= s_Energy_Bin_739;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_739 <= '0';
      end if;
    end if;
  end process  Energy_Bin_739;         
  
     Energy_Bin_740 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_740   <=  (others =>'0');
		Energy_Bin_Rdy_740 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E740_C1_L and PEAK_C1 <= s_E740_C1_H and Bin_OR = '0') then
         s_Energy_Bin_740 <= s_Energy_Bin_740 +'1';
		 Energy_Bin_Rdy_740 <= '1';
		else
		 s_Energy_Bin_740 <= s_Energy_Bin_740;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_740 <= '0';
      end if;
    end if;
  end process  Energy_Bin_740;    
  
  Energy_Bin_741 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_741   <=  (others =>'0');
		Energy_Bin_Rdy_741 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E741_C1_L and PEAK_C1 <= s_E741_C1_H and Bin_OR = '0') then
         s_Energy_Bin_741 <= s_Energy_Bin_741 +'1';
		 Energy_Bin_Rdy_741 <= '1';
		else
		 s_Energy_Bin_741 <= s_Energy_Bin_741;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_741 <= '0';
      end if;
    end if;
  end process  Energy_Bin_741;   
  
  Energy_Bin_742 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_742   <=  (others =>'0');
	    Energy_Bin_Rdy_742 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E742_C1_L and PEAK_C1 <= s_E742_C1_H and Bin_OR = '0') then
         s_Energy_Bin_742 <= s_Energy_Bin_742 +'1';
		 Energy_Bin_Rdy_742 <= '1';
		else
		 s_Energy_Bin_742 <= s_Energy_Bin_742;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_742 <= '0';
      end if;
    end if;
  end process  Energy_Bin_742;   
  
  Energy_Bin_743 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_743   <=  (others =>'0');
	    Energy_Bin_Rdy_743 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E743_C1_L and PEAK_C1 <= s_E743_C1_H and Bin_OR = '0') then
         s_Energy_Bin_743 <= s_Energy_Bin_743 +'1';
		 Energy_Bin_Rdy_743 <= '1';
		else
		 s_Energy_Bin_743 <= s_Energy_Bin_743;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_743 <= '0';
      end if;
    end if;
  end process  Energy_Bin_743;   
  
  Energy_Bin_744 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_744   <=  (others =>'0');
		Energy_Bin_Rdy_744 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E744_C1_L and PEAK_C1 <= s_E744_C1_H and Bin_OR = '0') then
         s_Energy_Bin_744 <= s_Energy_Bin_744 +'1';
		 Energy_Bin_Rdy_744 <= '1';
		else
		 s_Energy_Bin_744 <= s_Energy_Bin_744;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_744 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_744;   
 
 
  Energy_Bin_745 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_745   <=  (others =>'0');
		Energy_Bin_Rdy_745 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E745_C1_L and PEAK_C1 <= s_E745_C1_H and Bin_OR = '0') then
         s_Energy_Bin_745 <= s_Energy_Bin_745 +'1';
		 Energy_Bin_Rdy_745 <= '1';
		else
		 s_Energy_Bin_745 <= s_Energy_Bin_745;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_745 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_745;  
 
  
  Energy_Bin_746 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_746   <=  (others =>'0');
		Energy_Bin_Rdy_746 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E746_C1_L and PEAK_C1 <= s_E746_C1_H and Bin_OR = '0') then
         s_Energy_Bin_746 <= s_Energy_Bin_746 +'1';
		 Energy_Bin_Rdy_746 <= '1';
		else
		 s_Energy_Bin_746 <= s_Energy_Bin_746;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_746 <= '0';
      end if;
    end if;
  end process  Energy_Bin_746;   
  
 Energy_Bin_747 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_747   <=  (others =>'0');
		Energy_Bin_Rdy_747 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E747_C1_L and PEAK_C1 <= s_E747_C1_H and Bin_OR = '0') then
         s_Energy_Bin_747 <= s_Energy_Bin_747 +'1';
		 Energy_Bin_Rdy_747 <= '1';
		else
		 s_Energy_Bin_747 <= s_Energy_Bin_747;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_747 <= '0';
      end if;
    end if;
  end process  Energy_Bin_747;   
  
  Energy_Bin_748 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_748   <=  (others =>'0');
		Energy_Bin_Rdy_748 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E748_C1_L and PEAK_C1 <= s_E748_C1_H and Bin_OR = '0') then
         s_Energy_Bin_748 <= s_Energy_Bin_748 +'1';
		 Energy_Bin_Rdy_748 <= '1';
		else
		 s_Energy_Bin_748 <= s_Energy_Bin_748;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_748 <= '0';
      end if;
    end if;
  end process  Energy_Bin_748;   
  
  Energy_Bin_749 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_749   <=  (others =>'0');
		Energy_Bin_Rdy_749 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E749_C1_L and PEAK_C1 <= s_E749_C1_H and Bin_OR = '0') then
         s_Energy_Bin_749 <= s_Energy_Bin_749 +'1';
		 Energy_Bin_Rdy_749 <= '1';
		else
		 s_Energy_Bin_749 <= s_Energy_Bin_749;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_749 <= '0';
      end if;
    end if;
  end process  Energy_Bin_749;          
  
  
     Energy_Bin_750 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_750   <=  (others =>'0');
		Energy_Bin_Rdy_750 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E750_C1_L and PEAK_C1 <= s_E750_C1_H and Bin_OR = '0') then
         s_Energy_Bin_750 <= s_Energy_Bin_750 +'1';
		 Energy_Bin_Rdy_750 <= '1';
		else
		 s_Energy_Bin_750 <= s_Energy_Bin_750;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_750 <= '0';
      end if;
    end if;
  end process  Energy_Bin_750;    
  
  Energy_Bin_751 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_751   <=  (others =>'0');
		Energy_Bin_Rdy_751 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E751_C1_L and PEAK_C1 <= s_E751_C1_H and Bin_OR = '0') then
         s_Energy_Bin_751 <= s_Energy_Bin_751 +'1';
		 Energy_Bin_Rdy_751 <= '1';
		else
		 s_Energy_Bin_751 <= s_Energy_Bin_751;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_751 <= '0';
      end if;
    end if;
  end process  Energy_Bin_751;   
  
  Energy_Bin_752 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_752   <=  (others =>'0');
	    Energy_Bin_Rdy_752 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E752_C1_L and PEAK_C1 <= s_E752_C1_H and Bin_OR = '0') then
         s_Energy_Bin_752 <= s_Energy_Bin_752 +'1';
		 Energy_Bin_Rdy_752 <= '1';
		else
		 s_Energy_Bin_752 <= s_Energy_Bin_752;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_752 <= '0';
      end if;
    end if;
  end process  Energy_Bin_752;   
  
  Energy_Bin_753 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_753   <=  (others =>'0');
	    Energy_Bin_Rdy_753 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E753_C1_L and PEAK_C1 <= s_E753_C1_H and Bin_OR = '0') then
         s_Energy_Bin_753 <= s_Energy_Bin_753 +'1';
		 Energy_Bin_Rdy_753 <= '1';
		else
		 s_Energy_Bin_753 <= s_Energy_Bin_753;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_753 <= '0';
      end if;
    end if;
  end process  Energy_Bin_753;   
  
  Energy_Bin_754 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_754   <=  (others =>'0');
		Energy_Bin_Rdy_754 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E754_C1_L and PEAK_C1 <= s_E754_C1_H and Bin_OR = '0') then
         s_Energy_Bin_754 <= s_Energy_Bin_754 +'1';
		 Energy_Bin_Rdy_754 <= '1';
		else
		 s_Energy_Bin_754 <= s_Energy_Bin_754;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_754 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_754;   
 
 
  Energy_Bin_755 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_755   <=  (others =>'0');
		Energy_Bin_Rdy_755 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E755_C1_L and PEAK_C1 <= s_E755_C1_H and Bin_OR = '0') then
         s_Energy_Bin_755 <= s_Energy_Bin_755 +'1';
		 Energy_Bin_Rdy_755 <= '1';
		else
		 s_Energy_Bin_755 <= s_Energy_Bin_755;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_755 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_755;  
 
  
  Energy_Bin_756 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_756   <=  (others =>'0');
		Energy_Bin_Rdy_756 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E756_C1_L and PEAK_C1 <= s_E756_C1_H and Bin_OR = '0') then
         s_Energy_Bin_756 <= s_Energy_Bin_756 +'1';
		 Energy_Bin_Rdy_756 <= '1';
		else
		 s_Energy_Bin_756 <= s_Energy_Bin_756;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_756 <= '0';
      end if;
    end if;
  end process  Energy_Bin_756;   
  
 Energy_Bin_757 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_757   <=  (others =>'0');
		Energy_Bin_Rdy_757 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E757_C1_L and PEAK_C1 <= s_E757_C1_H and Bin_OR = '0') then
         s_Energy_Bin_757 <= s_Energy_Bin_757 +'1';
		 Energy_Bin_Rdy_757 <= '1';
		else
		 s_Energy_Bin_757 <= s_Energy_Bin_757;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_757 <= '0';
      end if;
    end if;
  end process  Energy_Bin_757;   
  
  Energy_Bin_758 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_758   <=  (others =>'0');
		Energy_Bin_Rdy_758 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E758_C1_L and PEAK_C1 <= s_E758_C1_H and Bin_OR = '0') then
         s_Energy_Bin_758 <= s_Energy_Bin_758 +'1';
		 Energy_Bin_Rdy_758 <= '1';
		else
		 s_Energy_Bin_758 <= s_Energy_Bin_758;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_758 <= '0';
      end if;
    end if;
  end process  Energy_Bin_758;   
  
  Energy_Bin_759 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_759   <=  (others =>'0');
		Energy_Bin_Rdy_759 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E759_C1_L and PEAK_C1 <= s_E759_C1_H and Bin_OR = '0') then
         s_Energy_Bin_759 <= s_Energy_Bin_759 +'1';
		 Energy_Bin_Rdy_759 <= '1';
		else
		 s_Energy_Bin_759 <= s_Energy_Bin_759;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_759 <= '0';
      end if;
    end if;
  end process  Energy_Bin_759;           
  
     Energy_Bin_760 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_760   <=  (others =>'0');
		Energy_Bin_Rdy_760 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E760_C1_L and PEAK_C1 <= s_E760_C1_H and Bin_OR = '0') then
         s_Energy_Bin_760 <= s_Energy_Bin_760 +'1';
		 Energy_Bin_Rdy_760 <= '1';
		else
		 s_Energy_Bin_760 <= s_Energy_Bin_760;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_760 <= '0';
      end if;
    end if;
  end process  Energy_Bin_760;    
  
  Energy_Bin_761 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_761   <=  (others =>'0');
		Energy_Bin_Rdy_761 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E761_C1_L and PEAK_C1 <= s_E761_C1_H and Bin_OR = '0') then
         s_Energy_Bin_761 <= s_Energy_Bin_761 +'1';
		 Energy_Bin_Rdy_761 <= '1';
		else
		 s_Energy_Bin_761 <= s_Energy_Bin_761;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_761 <= '0';
      end if;
    end if;
  end process  Energy_Bin_761;   
  
  Energy_Bin_762 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_762   <=  (others =>'0');
	    Energy_Bin_Rdy_762 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E762_C1_L and PEAK_C1 <= s_E762_C1_H and Bin_OR = '0') then
         s_Energy_Bin_762 <= s_Energy_Bin_762 +'1';
		 Energy_Bin_Rdy_762 <= '1';
		else
		 s_Energy_Bin_762 <= s_Energy_Bin_762;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_762 <= '0';
      end if;
    end if;
  end process  Energy_Bin_762;   
  
  Energy_Bin_763 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_763   <=  (others =>'0');
	    Energy_Bin_Rdy_763 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E763_C1_L and PEAK_C1 <= s_E763_C1_H and Bin_OR = '0') then
         s_Energy_Bin_763 <= s_Energy_Bin_763 +'1';
		 Energy_Bin_Rdy_763 <= '1';
		else
		 s_Energy_Bin_763 <= s_Energy_Bin_763;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_763 <= '0';
      end if;
    end if;
  end process  Energy_Bin_763;   
  
  Energy_Bin_764 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_764   <=  (others =>'0');
		Energy_Bin_Rdy_764 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E764_C1_L and PEAK_C1 <= s_E764_C1_H and Bin_OR = '0') then
         s_Energy_Bin_764 <= s_Energy_Bin_764 +'1';
		 Energy_Bin_Rdy_764 <= '1';
		else
		 s_Energy_Bin_764 <= s_Energy_Bin_764;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_764 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_764;   
 
 
  Energy_Bin_765 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_765   <=  (others =>'0');
		Energy_Bin_Rdy_765 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E765_C1_L and PEAK_C1 <= s_E765_C1_H and Bin_OR = '0') then
         s_Energy_Bin_765 <= s_Energy_Bin_765 +'1';
		 Energy_Bin_Rdy_765 <= '1';
		else
		 s_Energy_Bin_765 <= s_Energy_Bin_765;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_765 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_765;  
 
  
  Energy_Bin_766 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_766   <=  (others =>'0');
		Energy_Bin_Rdy_766 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E766_C1_L and PEAK_C1 <= s_E766_C1_H and Bin_OR = '0') then
         s_Energy_Bin_766 <= s_Energy_Bin_766 +'1';
		 Energy_Bin_Rdy_766 <= '1';
		else
		 s_Energy_Bin_766 <= s_Energy_Bin_766;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_766 <= '0';
      end if;
    end if;
  end process  Energy_Bin_766;   
  
 Energy_Bin_767 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_767   <=  (others =>'0');
		Energy_Bin_Rdy_767 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E767_C1_L and PEAK_C1 <= s_E767_C1_H and Bin_OR = '0') then
         s_Energy_Bin_767 <= s_Energy_Bin_767 +'1';
		 Energy_Bin_Rdy_767 <= '1';
		else
		 s_Energy_Bin_767 <= s_Energy_Bin_767;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_767 <= '0';
      end if;
    end if;
  end process  Energy_Bin_767;   
  
  Energy_Bin_768 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_768   <=  (others =>'0');
		Energy_Bin_Rdy_768 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E768_C1_L and PEAK_C1 <= s_E768_C1_H and Bin_OR = '0') then
         s_Energy_Bin_768 <= s_Energy_Bin_768 +'1';
		 Energy_Bin_Rdy_768 <= '1';
		else
		 s_Energy_Bin_768 <= s_Energy_Bin_768;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_768 <= '0';
      end if;
    end if;
  end process  Energy_Bin_768;   
  
  Energy_Bin_769 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_769   <=  (others =>'0');
		Energy_Bin_Rdy_769 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E769_C1_L and PEAK_C1 <= s_E769_C1_H and Bin_OR = '0') then
         s_Energy_Bin_769 <= s_Energy_Bin_769 +'1';
		 Energy_Bin_Rdy_769 <= '1';
		else
		 s_Energy_Bin_769 <= s_Energy_Bin_769;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_769 <= '0';
      end if;
    end if;
  end process  Energy_Bin_769;         
  
     Energy_Bin_770 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_770   <=  (others =>'0');
		Energy_Bin_Rdy_770 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E770_C1_L and PEAK_C1 <= s_E770_C1_H and Bin_OR = '0') then
         s_Energy_Bin_770 <= s_Energy_Bin_770 +'1';
		 Energy_Bin_Rdy_770 <= '1';
		else
		 s_Energy_Bin_770 <= s_Energy_Bin_770;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_770 <= '0';
      end if;
    end if;
  end process  Energy_Bin_770;    
  
  Energy_Bin_771 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_771   <=  (others =>'0');
		Energy_Bin_Rdy_771 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E771_C1_L and PEAK_C1 <= s_E771_C1_H and Bin_OR = '0') then
         s_Energy_Bin_771 <= s_Energy_Bin_771 +'1';
		 Energy_Bin_Rdy_771 <= '1';
		else
		 s_Energy_Bin_771 <= s_Energy_Bin_771;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_771 <= '0';
      end if;
    end if;
  end process  Energy_Bin_771;   
  
  Energy_Bin_772 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_772   <=  (others =>'0');
	    Energy_Bin_Rdy_772 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E772_C1_L and PEAK_C1 <= s_E772_C1_H and Bin_OR = '0') then
         s_Energy_Bin_772 <= s_Energy_Bin_772 +'1';
		 Energy_Bin_Rdy_772 <= '1';
		else
		 s_Energy_Bin_772 <= s_Energy_Bin_772;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_772 <= '0';
      end if;
    end if;
  end process  Energy_Bin_772;   
  
  Energy_Bin_773 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_773   <=  (others =>'0');
	    Energy_Bin_Rdy_773 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E773_C1_L and PEAK_C1 <= s_E773_C1_H and Bin_OR = '0') then
         s_Energy_Bin_773 <= s_Energy_Bin_773 +'1';
		 Energy_Bin_Rdy_773 <= '1';
		else
		 s_Energy_Bin_773 <= s_Energy_Bin_773;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_773 <= '0';
      end if;
    end if;
  end process  Energy_Bin_773;   
  
  Energy_Bin_774 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_774   <=  (others =>'0');
		Energy_Bin_Rdy_774 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E774_C1_L and PEAK_C1 <= s_E774_C1_H and Bin_OR = '0') then
         s_Energy_Bin_774 <= s_Energy_Bin_774 +'1';
		 Energy_Bin_Rdy_774 <= '1';
		else
		 s_Energy_Bin_774 <= s_Energy_Bin_774;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_774 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_774;   
 
 
  Energy_Bin_775 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_775   <=  (others =>'0');
		Energy_Bin_Rdy_775 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E775_C1_L and PEAK_C1 <= s_E775_C1_H and Bin_OR = '0') then
         s_Energy_Bin_775 <= s_Energy_Bin_775 +'1';
		 Energy_Bin_Rdy_775 <= '1';
		else
		 s_Energy_Bin_775 <= s_Energy_Bin_775;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_775 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_775;  
 
  
  Energy_Bin_776 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_776   <=  (others =>'0');
		Energy_Bin_Rdy_776 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E776_C1_L and PEAK_C1 <= s_E776_C1_H and Bin_OR = '0') then
         s_Energy_Bin_776 <= s_Energy_Bin_776 +'1';
		 Energy_Bin_Rdy_776 <= '1';
		else
		 s_Energy_Bin_776 <= s_Energy_Bin_776;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_776 <= '0';
      end if;
    end if;
  end process  Energy_Bin_776;   
  
 Energy_Bin_777 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_777   <=  (others =>'0');
		Energy_Bin_Rdy_777 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E777_C1_L and PEAK_C1 <= s_E777_C1_H and Bin_OR = '0') then
         s_Energy_Bin_777 <= s_Energy_Bin_777 +'1';
		 Energy_Bin_Rdy_777 <= '1';
		else
		 s_Energy_Bin_777 <= s_Energy_Bin_777;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_777 <= '0';
      end if;
    end if;
  end process  Energy_Bin_777;   
  
  Energy_Bin_778 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_778   <=  (others =>'0');
		Energy_Bin_Rdy_778 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E778_C1_L and PEAK_C1 <= s_E778_C1_H and Bin_OR = '0') then
         s_Energy_Bin_778 <= s_Energy_Bin_778 +'1';
		 Energy_Bin_Rdy_778 <= '1';
		else
		 s_Energy_Bin_778 <= s_Energy_Bin_778;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_778 <= '0';
      end if;
    end if;
  end process  Energy_Bin_778;   
  
  Energy_Bin_779 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_779   <=  (others =>'0');
		Energy_Bin_Rdy_779 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E779_C1_L and PEAK_C1 <= s_E779_C1_H and Bin_OR = '0') then
         s_Energy_Bin_779 <= s_Energy_Bin_779 +'1';
		 Energy_Bin_Rdy_779 <= '1';
		else
		 s_Energy_Bin_779 <= s_Energy_Bin_779;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_779 <= '0';
      end if;
    end if;
  end process  Energy_Bin_779;       
  
     Energy_Bin_780 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_780   <=  (others =>'0');
		Energy_Bin_Rdy_780 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E780_C1_L and PEAK_C1 <= s_E780_C1_H and Bin_OR = '0') then
         s_Energy_Bin_780 <= s_Energy_Bin_780 +'1';
		 Energy_Bin_Rdy_780 <= '1';
		else
		 s_Energy_Bin_780 <= s_Energy_Bin_780;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_780 <= '0';
      end if;
    end if;
  end process  Energy_Bin_780;    
  
  Energy_Bin_781 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_781   <=  (others =>'0');
		Energy_Bin_Rdy_781 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E781_C1_L and PEAK_C1 <= s_E781_C1_H and Bin_OR = '0') then
         s_Energy_Bin_781 <= s_Energy_Bin_781 +'1';
		 Energy_Bin_Rdy_781 <= '1';
		else
		 s_Energy_Bin_781 <= s_Energy_Bin_781;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_781 <= '0';
      end if;
    end if;
  end process  Energy_Bin_781;   
  
  Energy_Bin_782 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_782   <=  (others =>'0');
	    Energy_Bin_Rdy_782 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E782_C1_L and PEAK_C1 <= s_E782_C1_H and Bin_OR = '0') then
         s_Energy_Bin_782 <= s_Energy_Bin_782 +'1';
		 Energy_Bin_Rdy_782 <= '1';
		else
		 s_Energy_Bin_782 <= s_Energy_Bin_782;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_782 <= '0';
      end if;
    end if;
  end process  Energy_Bin_782;   
  
  Energy_Bin_783 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_783   <=  (others =>'0');
	    Energy_Bin_Rdy_783 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E783_C1_L and PEAK_C1 <= s_E783_C1_H and Bin_OR = '0') then
         s_Energy_Bin_783 <= s_Energy_Bin_783 +'1';
		 Energy_Bin_Rdy_783 <= '1';
		else
		 s_Energy_Bin_783 <= s_Energy_Bin_783;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_783 <= '0';
      end if;
    end if;
  end process  Energy_Bin_783;   
  
  Energy_Bin_784 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_784   <=  (others =>'0');
		Energy_Bin_Rdy_784 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E784_C1_L and PEAK_C1 <= s_E784_C1_H and Bin_OR = '0') then
         s_Energy_Bin_784 <= s_Energy_Bin_784 +'1';
		 Energy_Bin_Rdy_784 <= '1';
		else
		 s_Energy_Bin_784 <= s_Energy_Bin_784;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_784 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_784;   
 
 
  Energy_Bin_785 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_785   <=  (others =>'0');
		Energy_Bin_Rdy_785 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E785_C1_L and PEAK_C1 <= s_E785_C1_H and Bin_OR = '0') then
         s_Energy_Bin_785 <= s_Energy_Bin_785 +'1';
		 Energy_Bin_Rdy_785 <= '1';
		else
		 s_Energy_Bin_785 <= s_Energy_Bin_785;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_785 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_785;  
 
  
  Energy_Bin_786 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_786   <=  (others =>'0');
		Energy_Bin_Rdy_786 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E786_C1_L and PEAK_C1 <= s_E786_C1_H and Bin_OR = '0') then
         s_Energy_Bin_786 <= s_Energy_Bin_786 +'1';
		 Energy_Bin_Rdy_786 <= '1';
		else
		 s_Energy_Bin_786 <= s_Energy_Bin_786;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_786 <= '0';
      end if;
    end if;
  end process  Energy_Bin_786;   
  
 Energy_Bin_787 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_787   <=  (others =>'0');
		Energy_Bin_Rdy_787 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E787_C1_L and PEAK_C1 <= s_E787_C1_H and Bin_OR = '0') then
         s_Energy_Bin_787 <= s_Energy_Bin_787 +'1';
		 Energy_Bin_Rdy_787 <= '1';
		else
		 s_Energy_Bin_787 <= s_Energy_Bin_787;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_787 <= '0';
      end if;
    end if;
  end process  Energy_Bin_787;   
  
  Energy_Bin_788 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_788   <=  (others =>'0');
		Energy_Bin_Rdy_788 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E788_C1_L and PEAK_C1 <= s_E788_C1_H and Bin_OR = '0') then
         s_Energy_Bin_788 <= s_Energy_Bin_788 +'1';
		 Energy_Bin_Rdy_788 <= '1';
		else
		 s_Energy_Bin_788 <= s_Energy_Bin_788;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_788 <= '0';
      end if;
    end if;
  end process  Energy_Bin_788;   
  
  Energy_Bin_789 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_789   <=  (others =>'0');
		Energy_Bin_Rdy_789 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E789_C1_L and PEAK_C1 <= s_E789_C1_H and Bin_OR = '0') then
         s_Energy_Bin_789 <= s_Energy_Bin_789 +'1';
		 Energy_Bin_Rdy_789 <= '1';
		else
		 s_Energy_Bin_789 <= s_Energy_Bin_789;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_789 <= '0';
      end if;
    end if;
  end process  Energy_Bin_789;      
  
     Energy_Bin_790 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_790   <=  (others =>'0');
		Energy_Bin_Rdy_790 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E790_C1_L and PEAK_C1 <= s_E790_C1_H and Bin_OR = '0') then
         s_Energy_Bin_790 <= s_Energy_Bin_790 +'1';
		 Energy_Bin_Rdy_790 <= '1';
		else
		 s_Energy_Bin_790 <= s_Energy_Bin_790;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_790 <= '0';
      end if;
    end if;
  end process  Energy_Bin_790;    
  
  Energy_Bin_791 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_791   <=  (others =>'0');
		Energy_Bin_Rdy_791 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E791_C1_L and PEAK_C1 <= s_E791_C1_H and Bin_OR = '0') then
         s_Energy_Bin_791 <= s_Energy_Bin_791 +'1';
		 Energy_Bin_Rdy_791 <= '1';
		else
		 s_Energy_Bin_791 <= s_Energy_Bin_791;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_791 <= '0';
      end if;
    end if;
  end process  Energy_Bin_791;   
  
  Energy_Bin_792 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_792   <=  (others =>'0');
	    Energy_Bin_Rdy_792 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E792_C1_L and PEAK_C1 <= s_E792_C1_H and Bin_OR = '0') then
         s_Energy_Bin_792 <= s_Energy_Bin_792 +'1';
		 Energy_Bin_Rdy_792 <= '1';
		else
		 s_Energy_Bin_792 <= s_Energy_Bin_792;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_792 <= '0';
      end if;
    end if;
  end process  Energy_Bin_792;   
  
  Energy_Bin_793 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_793   <=  (others =>'0');
	    Energy_Bin_Rdy_793 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E793_C1_L and PEAK_C1 <= s_E793_C1_H and Bin_OR = '0') then
         s_Energy_Bin_793 <= s_Energy_Bin_793 +'1';
		 Energy_Bin_Rdy_793 <= '1';
		else
		 s_Energy_Bin_793 <= s_Energy_Bin_793;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_793 <= '0';
      end if;
    end if;
  end process  Energy_Bin_793;   
  
  Energy_Bin_794 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_794   <=  (others =>'0');
		Energy_Bin_Rdy_794 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E794_C1_L and PEAK_C1 <= s_E794_C1_H and Bin_OR = '0') then
         s_Energy_Bin_794 <= s_Energy_Bin_794 +'1';
		 Energy_Bin_Rdy_794 <= '1';
		else
		 s_Energy_Bin_794 <= s_Energy_Bin_794;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_794 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_794;   
 
 
  Energy_Bin_795 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_795   <=  (others =>'0');
		Energy_Bin_Rdy_795 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E795_C1_L and PEAK_C1 <= s_E795_C1_H and Bin_OR = '0') then
         s_Energy_Bin_795 <= s_Energy_Bin_795 +'1';
		 Energy_Bin_Rdy_795 <= '1';
		else
		 s_Energy_Bin_795 <= s_Energy_Bin_795;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_795 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_795;  
 
  
  Energy_Bin_796 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_796   <=  (others =>'0');
		Energy_Bin_Rdy_796 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E796_C1_L and PEAK_C1 <= s_E796_C1_H and Bin_OR = '0') then
         s_Energy_Bin_796 <= s_Energy_Bin_796 +'1';
		 Energy_Bin_Rdy_796 <= '1';
		else
		 s_Energy_Bin_796 <= s_Energy_Bin_796;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_796 <= '0';
      end if;
    end if;
  end process  Energy_Bin_796;   
  
 Energy_Bin_797 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_797   <=  (others =>'0');
		Energy_Bin_Rdy_797 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E797_C1_L and PEAK_C1 <= s_E797_C1_H and Bin_OR = '0') then
         s_Energy_Bin_797 <= s_Energy_Bin_797 +'1';
		 Energy_Bin_Rdy_797 <= '1';
		else
		 s_Energy_Bin_797 <= s_Energy_Bin_797;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_797 <= '0';
      end if;
    end if;
  end process  Energy_Bin_797;   
  
  Energy_Bin_798 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_798   <=  (others =>'0');
		Energy_Bin_Rdy_798 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E798_C1_L and PEAK_C1 <= s_E798_C1_H and Bin_OR = '0') then
         s_Energy_Bin_798 <= s_Energy_Bin_798 +'1';
		 Energy_Bin_Rdy_798 <= '1';
		else
		 s_Energy_Bin_798 <= s_Energy_Bin_798;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_798 <= '0';
      end if;
    end if;
  end process  Energy_Bin_798;   
  
  Energy_Bin_799 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_799   <=  (others =>'0');
		Energy_Bin_Rdy_799 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E799_C1_L and PEAK_C1 <= s_E799_C1_H and Bin_OR = '0') then
         s_Energy_Bin_799 <= s_Energy_Bin_799 +'1';
		 Energy_Bin_Rdy_799 <= '1';
		else
		 s_Energy_Bin_799 <= s_Energy_Bin_799;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_799 <= '0';
      end if;
    end if;
  end process  Energy_Bin_799;   

    Energy_Bin_800 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_800   <=  (others =>'0');
		Energy_Bin_Rdy_800 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E800_C1_L and PEAK_C1 <= s_E800_C1_H and Bin_OR = '0') then
         s_Energy_Bin_800 <= s_Energy_Bin_800 +'1';
		 Energy_Bin_Rdy_800 <= '1';
		else
		 s_Energy_Bin_800 <= s_Energy_Bin_800;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_800 <= '0';
      end if;
    end if;
  end process  Energy_Bin_800;    
  
  Energy_Bin_801 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_801   <=  (others =>'0');
		Energy_Bin_Rdy_801 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E801_C1_L and PEAK_C1 <= s_E801_C1_H and Bin_OR = '0') then
         s_Energy_Bin_801 <= s_Energy_Bin_801 +'1';
		 Energy_Bin_Rdy_801 <= '1';
		else
		 s_Energy_Bin_801 <= s_Energy_Bin_801;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_801 <= '0';
      end if;
    end if;
  end process  Energy_Bin_801;   
  
  Energy_Bin_802 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_802   <=  (others =>'0');
	    Energy_Bin_Rdy_802 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E802_C1_L and PEAK_C1 <= s_E802_C1_H and Bin_OR = '0') then
         s_Energy_Bin_802 <= s_Energy_Bin_802 +'1';
		 Energy_Bin_Rdy_802 <= '1';
		else
		 s_Energy_Bin_802 <= s_Energy_Bin_802;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_802 <= '0';
      end if;
    end if;
  end process  Energy_Bin_802;   
  
  Energy_Bin_803 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_803   <=  (others =>'0');
	    Energy_Bin_Rdy_803 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E803_C1_L and PEAK_C1 <= s_E803_C1_H and Bin_OR = '0') then
         s_Energy_Bin_803 <= s_Energy_Bin_803 +'1';
		 Energy_Bin_Rdy_803 <= '1';
		else
		 s_Energy_Bin_803 <= s_Energy_Bin_803;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_803 <= '0';
      end if;
    end if;
  end process  Energy_Bin_803;   
  
  Energy_Bin_804 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_804   <=  (others =>'0');
		Energy_Bin_Rdy_804 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E804_C1_L and PEAK_C1 <= s_E804_C1_H and Bin_OR = '0') then
         s_Energy_Bin_804 <= s_Energy_Bin_804 +'1';
		 Energy_Bin_Rdy_804 <= '1';
		else
		 s_Energy_Bin_804 <= s_Energy_Bin_804;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_804 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_804;   
 
 
  Energy_Bin_805 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_805   <=  (others =>'0');
		Energy_Bin_Rdy_805 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E805_C1_L and PEAK_C1 <= s_E805_C1_H and Bin_OR = '0') then
         s_Energy_Bin_805 <= s_Energy_Bin_805 +'1';
		 Energy_Bin_Rdy_805 <= '1';
		else
		 s_Energy_Bin_805 <= s_Energy_Bin_805;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_805 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_805;  
 
  
  Energy_Bin_806 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_806   <=  (others =>'0');
		Energy_Bin_Rdy_806 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E806_C1_L and PEAK_C1 <= s_E806_C1_H and Bin_OR = '0') then
         s_Energy_Bin_806 <= s_Energy_Bin_806 +'1';
		 Energy_Bin_Rdy_806 <= '1';
		else
		 s_Energy_Bin_806 <= s_Energy_Bin_806;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_806 <= '0';
      end if;
    end if;
  end process  Energy_Bin_806;   
  
 Energy_Bin_807 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_807   <=  (others =>'0');
		Energy_Bin_Rdy_807 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E807_C1_L and PEAK_C1 <= s_E807_C1_H and Bin_OR = '0') then
         s_Energy_Bin_807 <= s_Energy_Bin_807 +'1';
		 Energy_Bin_Rdy_807 <= '1';
		else
		 s_Energy_Bin_807 <= s_Energy_Bin_807;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_807 <= '0';
      end if;
    end if;
  end process  Energy_Bin_807;   
  
  Energy_Bin_808 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_808   <=  (others =>'0');
		Energy_Bin_Rdy_808 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E808_C1_L and PEAK_C1 <= s_E808_C1_H and Bin_OR = '0') then
         s_Energy_Bin_808 <= s_Energy_Bin_808 +'1';
		 Energy_Bin_Rdy_808 <= '1';
		else
		 s_Energy_Bin_808 <= s_Energy_Bin_808;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_808 <= '0';
      end if;
    end if;
  end process  Energy_Bin_808;   
  
  Energy_Bin_809 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_809   <=  (others =>'0');
		Energy_Bin_Rdy_809 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E809_C1_L and PEAK_C1 <= s_E809_C1_H and Bin_OR = '0') then
         s_Energy_Bin_809 <= s_Energy_Bin_809 +'1';
		 Energy_Bin_Rdy_809 <= '1';
		else
		 s_Energy_Bin_809 <= s_Energy_Bin_809;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_809 <= '0';
      end if;
    end if;
  end process  Energy_Bin_809;      
  
     Energy_Bin_810 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_810   <=  (others =>'0');
		Energy_Bin_Rdy_810 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E810_C1_L and PEAK_C1 <= s_E810_C1_H and Bin_OR = '0') then
         s_Energy_Bin_810 <= s_Energy_Bin_810 +'1';
		 Energy_Bin_Rdy_810 <= '1';
		else
		 s_Energy_Bin_810 <= s_Energy_Bin_810;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_810 <= '0';
      end if;
    end if;
  end process  Energy_Bin_810;    
  
  Energy_Bin_811 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_811   <=  (others =>'0');
		Energy_Bin_Rdy_811 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E811_C1_L and PEAK_C1 <= s_E811_C1_H and Bin_OR = '0') then
         s_Energy_Bin_811 <= s_Energy_Bin_811 +'1';
		 Energy_Bin_Rdy_811 <= '1';
		else
		 s_Energy_Bin_811 <= s_Energy_Bin_811;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_811 <= '0';
      end if;
    end if;
  end process  Energy_Bin_811;   
  
  Energy_Bin_812 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_812   <=  (others =>'0');
	    Energy_Bin_Rdy_812 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E812_C1_L and PEAK_C1 <= s_E812_C1_H and Bin_OR = '0') then
         s_Energy_Bin_812 <= s_Energy_Bin_812 +'1';
		 Energy_Bin_Rdy_812 <= '1';
		else
		 s_Energy_Bin_812 <= s_Energy_Bin_812;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_812 <= '0';
      end if;
    end if;
  end process  Energy_Bin_812;   
  
  Energy_Bin_813 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_813   <=  (others =>'0');
	    Energy_Bin_Rdy_813 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E813_C1_L and PEAK_C1 <= s_E813_C1_H and Bin_OR = '0') then
         s_Energy_Bin_813 <= s_Energy_Bin_813 +'1';
		 Energy_Bin_Rdy_813 <= '1';
		else
		 s_Energy_Bin_813 <= s_Energy_Bin_813;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_813 <= '0';
      end if;
    end if;
  end process  Energy_Bin_813;   
  
  Energy_Bin_814 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_814   <=  (others =>'0');
		Energy_Bin_Rdy_814 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E814_C1_L and PEAK_C1 <= s_E814_C1_H and Bin_OR = '0') then
         s_Energy_Bin_814 <= s_Energy_Bin_814 +'1';
		 Energy_Bin_Rdy_814 <= '1';
		else
		 s_Energy_Bin_814 <= s_Energy_Bin_814;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_814 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_814;   
 
 
  Energy_Bin_815 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_815   <=  (others =>'0');
		Energy_Bin_Rdy_815 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E815_C1_L and PEAK_C1 <= s_E815_C1_H and Bin_OR = '0') then
         s_Energy_Bin_815 <= s_Energy_Bin_815 +'1';
		 Energy_Bin_Rdy_815 <= '1';
		else
		 s_Energy_Bin_815 <= s_Energy_Bin_815;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_815 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_815;  
 
  
  Energy_Bin_816 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_816   <=  (others =>'0');
		Energy_Bin_Rdy_816 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E816_C1_L and PEAK_C1 <= s_E816_C1_H and Bin_OR = '0') then
         s_Energy_Bin_816 <= s_Energy_Bin_816 +'1';
		 Energy_Bin_Rdy_816 <= '1';
		else
		 s_Energy_Bin_816 <= s_Energy_Bin_816;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_816 <= '0';
      end if;
    end if;
  end process  Energy_Bin_816;   
  
 Energy_Bin_817 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_817   <=  (others =>'0');
		Energy_Bin_Rdy_817 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E817_C1_L and PEAK_C1 <= s_E817_C1_H and Bin_OR = '0') then
         s_Energy_Bin_817 <= s_Energy_Bin_817 +'1';
		 Energy_Bin_Rdy_817 <= '1';
		else
		 s_Energy_Bin_817 <= s_Energy_Bin_817;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_817 <= '0';
      end if;
    end if;
  end process  Energy_Bin_817;   
  
  Energy_Bin_818 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_818   <=  (others =>'0');
		Energy_Bin_Rdy_818 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E818_C1_L and PEAK_C1 <= s_E818_C1_H and Bin_OR = '0') then
         s_Energy_Bin_818 <= s_Energy_Bin_818 +'1';
		 Energy_Bin_Rdy_818 <= '1';
		else
		 s_Energy_Bin_818 <= s_Energy_Bin_818;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_818 <= '0';
      end if;
    end if;
  end process  Energy_Bin_818;   
  
  Energy_Bin_819 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_819   <=  (others =>'0');
		Energy_Bin_Rdy_819 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E819_C1_L and PEAK_C1 <= s_E819_C1_H and Bin_OR = '0') then
         s_Energy_Bin_819 <= s_Energy_Bin_819 +'1';
		 Energy_Bin_Rdy_819 <= '1';
		else
		 s_Energy_Bin_819 <= s_Energy_Bin_819;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_819 <= '0';
      end if;
    end if;
  end process  Energy_Bin_819;       
  
     Energy_Bin_820 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_820   <=  (others =>'0');
		Energy_Bin_Rdy_820 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E820_C1_L and PEAK_C1 <= s_E820_C1_H and Bin_OR = '0') then
         s_Energy_Bin_820 <= s_Energy_Bin_820 +'1';
		 Energy_Bin_Rdy_820 <= '1';
		else
		 s_Energy_Bin_820 <= s_Energy_Bin_820;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_820 <= '0';
      end if;
    end if;
  end process  Energy_Bin_820;    
  
  Energy_Bin_821 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_821   <=  (others =>'0');
		Energy_Bin_Rdy_821 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E821_C1_L and PEAK_C1 <= s_E821_C1_H and Bin_OR = '0') then
         s_Energy_Bin_821 <= s_Energy_Bin_821 +'1';
		 Energy_Bin_Rdy_821 <= '1';
		else
		 s_Energy_Bin_821 <= s_Energy_Bin_821;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_821 <= '0';
      end if;
    end if;
  end process  Energy_Bin_821;   
  
  Energy_Bin_822 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_822   <=  (others =>'0');
	    Energy_Bin_Rdy_822 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E822_C1_L and PEAK_C1 <= s_E822_C1_H and Bin_OR = '0') then
         s_Energy_Bin_822 <= s_Energy_Bin_822 +'1';
		 Energy_Bin_Rdy_822 <= '1';
		else
		 s_Energy_Bin_822 <= s_Energy_Bin_822;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_822 <= '0';
      end if;
    end if;
  end process  Energy_Bin_822;   
  
  Energy_Bin_823 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_823   <=  (others =>'0');
	    Energy_Bin_Rdy_823 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E823_C1_L and PEAK_C1 <= s_E823_C1_H and Bin_OR = '0') then
         s_Energy_Bin_823 <= s_Energy_Bin_823 +'1';
		 Energy_Bin_Rdy_823 <= '1';
		else
		 s_Energy_Bin_823 <= s_Energy_Bin_823;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_823 <= '0';
      end if;
    end if;
  end process  Energy_Bin_823;   
  
  Energy_Bin_824 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_824   <=  (others =>'0');
		Energy_Bin_Rdy_824 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E824_C1_L and PEAK_C1 <= s_E824_C1_H and Bin_OR = '0') then
         s_Energy_Bin_824 <= s_Energy_Bin_824 +'1';
		 Energy_Bin_Rdy_824 <= '1';
		else
		 s_Energy_Bin_824 <= s_Energy_Bin_824;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_824 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_824;   
 
 
  Energy_Bin_825 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_825   <=  (others =>'0');
		Energy_Bin_Rdy_825 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E825_C1_L and PEAK_C1 <= s_E825_C1_H and Bin_OR = '0') then
         s_Energy_Bin_825 <= s_Energy_Bin_825 +'1';
		 Energy_Bin_Rdy_825 <= '1';
		else
		 s_Energy_Bin_825 <= s_Energy_Bin_825;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_825 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_825;  
 
  
  Energy_Bin_826 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_826   <=  (others =>'0');
		Energy_Bin_Rdy_826 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E826_C1_L and PEAK_C1 <= s_E826_C1_H and Bin_OR = '0') then
         s_Energy_Bin_826 <= s_Energy_Bin_826 +'1';
		 Energy_Bin_Rdy_826 <= '1';
		else
		 s_Energy_Bin_826 <= s_Energy_Bin_826;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_826 <= '0';
      end if;
    end if;
  end process  Energy_Bin_826;   
  
 Energy_Bin_827 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_827   <=  (others =>'0');
		Energy_Bin_Rdy_827 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E827_C1_L and PEAK_C1 <= s_E827_C1_H and Bin_OR = '0') then
         s_Energy_Bin_827 <= s_Energy_Bin_827 +'1';
		 Energy_Bin_Rdy_827 <= '1';
		else
		 s_Energy_Bin_827 <= s_Energy_Bin_827;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_827 <= '0';
      end if;
    end if;
  end process  Energy_Bin_827;   
  
  Energy_Bin_828 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_828   <=  (others =>'0');
		Energy_Bin_Rdy_828 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E828_C1_L and PEAK_C1 <= s_E828_C1_H and Bin_OR = '0') then
         s_Energy_Bin_828 <= s_Energy_Bin_828 +'1';
		 Energy_Bin_Rdy_828 <= '1';
		else
		 s_Energy_Bin_828 <= s_Energy_Bin_828;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_828 <= '0';
      end if;
    end if;
  end process  Energy_Bin_828;   
  
  Energy_Bin_829 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_829   <=  (others =>'0');
		Energy_Bin_Rdy_829 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E829_C1_L and PEAK_C1 <= s_E829_C1_H and Bin_OR = '0') then
         s_Energy_Bin_829 <= s_Energy_Bin_829 +'1';
		 Energy_Bin_Rdy_829 <= '1';
		else
		 s_Energy_Bin_829 <= s_Energy_Bin_829;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_829 <= '0';
      end if;
    end if;
  end process  Energy_Bin_829;        
  
     Energy_Bin_830 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_830   <=  (others =>'0');
		Energy_Bin_Rdy_830 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E830_C1_L and PEAK_C1 <= s_E830_C1_H and Bin_OR = '0') then
         s_Energy_Bin_830 <= s_Energy_Bin_830 +'1';
		 Energy_Bin_Rdy_830 <= '1';
		else
		 s_Energy_Bin_830 <= s_Energy_Bin_830;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_830 <= '0';
      end if;
    end if;
  end process  Energy_Bin_830;    
  
  Energy_Bin_831 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_831   <=  (others =>'0');
		Energy_Bin_Rdy_831 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E831_C1_L and PEAK_C1 <= s_E831_C1_H and Bin_OR = '0') then
         s_Energy_Bin_831 <= s_Energy_Bin_831 +'1';
		 Energy_Bin_Rdy_831 <= '1';
		else
		 s_Energy_Bin_831 <= s_Energy_Bin_831;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_831 <= '0';
      end if;
    end if;
  end process  Energy_Bin_831;   
  
  Energy_Bin_832 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_832   <=  (others =>'0');
	    Energy_Bin_Rdy_832 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E832_C1_L and PEAK_C1 <= s_E832_C1_H and Bin_OR = '0') then
         s_Energy_Bin_832 <= s_Energy_Bin_832 +'1';
		 Energy_Bin_Rdy_832 <= '1';
		else
		 s_Energy_Bin_832 <= s_Energy_Bin_832;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_832 <= '0';
      end if;
    end if;
  end process  Energy_Bin_832;   
  
  Energy_Bin_833 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_833   <=  (others =>'0');
	    Energy_Bin_Rdy_833 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E833_C1_L and PEAK_C1 <= s_E833_C1_H and Bin_OR = '0') then
         s_Energy_Bin_833 <= s_Energy_Bin_833 +'1';
		 Energy_Bin_Rdy_833 <= '1';
		else
		 s_Energy_Bin_833 <= s_Energy_Bin_833;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_833 <= '0';
      end if;
    end if;
  end process  Energy_Bin_833;   
  
  Energy_Bin_834 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_834   <=  (others =>'0');
		Energy_Bin_Rdy_834 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E834_C1_L and PEAK_C1 <= s_E834_C1_H and Bin_OR = '0') then
         s_Energy_Bin_834 <= s_Energy_Bin_834 +'1';
		 Energy_Bin_Rdy_834 <= '1';
		else
		 s_Energy_Bin_834 <= s_Energy_Bin_834;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_834 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_834;   
 
 
  Energy_Bin_835 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_835   <=  (others =>'0');
		Energy_Bin_Rdy_835 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E835_C1_L and PEAK_C1 <= s_E835_C1_H and Bin_OR = '0') then
         s_Energy_Bin_835 <= s_Energy_Bin_835 +'1';
		 Energy_Bin_Rdy_835 <= '1';
		else
		 s_Energy_Bin_835 <= s_Energy_Bin_835;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_835 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_835;  
 
  
  Energy_Bin_836 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_836   <=  (others =>'0');
		Energy_Bin_Rdy_836 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E836_C1_L and PEAK_C1 <= s_E836_C1_H and Bin_OR = '0') then
         s_Energy_Bin_836 <= s_Energy_Bin_836 +'1';
		 Energy_Bin_Rdy_836 <= '1';
		else
		 s_Energy_Bin_836 <= s_Energy_Bin_836;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_836 <= '0';
      end if;
    end if;
  end process  Energy_Bin_836;   
  
 Energy_Bin_837 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_837   <=  (others =>'0');
		Energy_Bin_Rdy_837 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E837_C1_L and PEAK_C1 <= s_E837_C1_H and Bin_OR = '0') then
         s_Energy_Bin_837 <= s_Energy_Bin_837 +'1';
		 Energy_Bin_Rdy_837 <= '1';
		else
		 s_Energy_Bin_837 <= s_Energy_Bin_837;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_837 <= '0';
      end if;
    end if;
  end process  Energy_Bin_837;   
  
  Energy_Bin_838 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_838   <=  (others =>'0');
		Energy_Bin_Rdy_838 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E838_C1_L and PEAK_C1 <= s_E838_C1_H and Bin_OR = '0') then
         s_Energy_Bin_838 <= s_Energy_Bin_838 +'1';
		 Energy_Bin_Rdy_838 <= '1';
		else
		 s_Energy_Bin_838 <= s_Energy_Bin_838;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_838 <= '0';
      end if;
    end if;
  end process  Energy_Bin_838;   
  
  Energy_Bin_839 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_839   <=  (others =>'0');
		Energy_Bin_Rdy_839 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E839_C1_L and PEAK_C1 <= s_E839_C1_H and Bin_OR = '0') then
         s_Energy_Bin_839 <= s_Energy_Bin_839 +'1';
		 Energy_Bin_Rdy_839 <= '1';
		else
		 s_Energy_Bin_839 <= s_Energy_Bin_839;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_839 <= '0';
      end if;
    end if;
  end process  Energy_Bin_839;         
  
     Energy_Bin_840 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_840   <=  (others =>'0');
		Energy_Bin_Rdy_840 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E840_C1_L and PEAK_C1 <= s_E840_C1_H and Bin_OR = '0') then
         s_Energy_Bin_840 <= s_Energy_Bin_840 +'1';
		 Energy_Bin_Rdy_840 <= '1';
		else
		 s_Energy_Bin_840 <= s_Energy_Bin_840;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_840 <= '0';
      end if;
    end if;
  end process  Energy_Bin_840;    
  
  Energy_Bin_841 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_841   <=  (others =>'0');
		Energy_Bin_Rdy_841 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E841_C1_L and PEAK_C1 <= s_E841_C1_H and Bin_OR = '0') then
         s_Energy_Bin_841 <= s_Energy_Bin_841 +'1';
		 Energy_Bin_Rdy_841 <= '1';
		else
		 s_Energy_Bin_841 <= s_Energy_Bin_841;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_841 <= '0';
      end if;
    end if;
  end process  Energy_Bin_841;   
  
  Energy_Bin_842 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_842   <=  (others =>'0');
	    Energy_Bin_Rdy_842 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E842_C1_L and PEAK_C1 <= s_E842_C1_H and Bin_OR = '0') then
         s_Energy_Bin_842 <= s_Energy_Bin_842 +'1';
		 Energy_Bin_Rdy_842 <= '1';
		else
		 s_Energy_Bin_842 <= s_Energy_Bin_842;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_842 <= '0';
      end if;
    end if;
  end process  Energy_Bin_842;   
  
  Energy_Bin_843 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_843   <=  (others =>'0');
	    Energy_Bin_Rdy_843 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E843_C1_L and PEAK_C1 <= s_E843_C1_H and Bin_OR = '0') then
         s_Energy_Bin_843 <= s_Energy_Bin_843 +'1';
		 Energy_Bin_Rdy_843 <= '1';
		else
		 s_Energy_Bin_843 <= s_Energy_Bin_843;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_843 <= '0';
      end if;
    end if;
  end process  Energy_Bin_843;   
  
  Energy_Bin_844 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_844   <=  (others =>'0');
		Energy_Bin_Rdy_844 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E844_C1_L and PEAK_C1 <= s_E844_C1_H and Bin_OR = '0') then
         s_Energy_Bin_844 <= s_Energy_Bin_844 +'1';
		 Energy_Bin_Rdy_844 <= '1';
		else
		 s_Energy_Bin_844 <= s_Energy_Bin_844;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_844 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_844;   
 
 
  Energy_Bin_845 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_845   <=  (others =>'0');
		Energy_Bin_Rdy_845 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E845_C1_L and PEAK_C1 <= s_E845_C1_H and Bin_OR = '0') then
         s_Energy_Bin_845 <= s_Energy_Bin_845 +'1';
		 Energy_Bin_Rdy_845 <= '1';
		else
		 s_Energy_Bin_845 <= s_Energy_Bin_845;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_845 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_845;  
 
  
  Energy_Bin_846 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_846   <=  (others =>'0');
		Energy_Bin_Rdy_846 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E846_C1_L and PEAK_C1 <= s_E846_C1_H and Bin_OR = '0') then
         s_Energy_Bin_846 <= s_Energy_Bin_846 +'1';
		 Energy_Bin_Rdy_846 <= '1';
		else
		 s_Energy_Bin_846 <= s_Energy_Bin_846;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_846 <= '0';
      end if;
    end if;
  end process  Energy_Bin_846;   
  
 Energy_Bin_847 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_847   <=  (others =>'0');
		Energy_Bin_Rdy_847 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E847_C1_L and PEAK_C1 <= s_E847_C1_H and Bin_OR = '0') then
         s_Energy_Bin_847 <= s_Energy_Bin_847 +'1';
		 Energy_Bin_Rdy_847 <= '1';
		else
		 s_Energy_Bin_847 <= s_Energy_Bin_847;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_847 <= '0';
      end if;
    end if;
  end process  Energy_Bin_847;   
  
  Energy_Bin_848 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_848   <=  (others =>'0');
		Energy_Bin_Rdy_848 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E848_C1_L and PEAK_C1 <= s_E848_C1_H and Bin_OR = '0') then
         s_Energy_Bin_848 <= s_Energy_Bin_848 +'1';
		 Energy_Bin_Rdy_848 <= '1';
		else
		 s_Energy_Bin_848 <= s_Energy_Bin_848;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_848 <= '0';
      end if;
    end if;
  end process  Energy_Bin_848;   
  
  Energy_Bin_849 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_849   <=  (others =>'0');
		Energy_Bin_Rdy_849 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E849_C1_L and PEAK_C1 <= s_E849_C1_H and Bin_OR = '0') then
         s_Energy_Bin_849 <= s_Energy_Bin_849 +'1';
		 Energy_Bin_Rdy_849 <= '1';
		else
		 s_Energy_Bin_849 <= s_Energy_Bin_849;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_849 <= '0';
      end if;
    end if;
  end process  Energy_Bin_849;          
  
  
     Energy_Bin_850 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_850   <=  (others =>'0');
		Energy_Bin_Rdy_850 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E850_C1_L and PEAK_C1 <= s_E850_C1_H and Bin_OR = '0') then
         s_Energy_Bin_850 <= s_Energy_Bin_850 +'1';
		 Energy_Bin_Rdy_850 <= '1';
		else
		 s_Energy_Bin_850 <= s_Energy_Bin_850;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_850 <= '0';
      end if;
    end if;
  end process  Energy_Bin_850;    
  
  Energy_Bin_851 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_851   <=  (others =>'0');
		Energy_Bin_Rdy_851 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E851_C1_L and PEAK_C1 <= s_E851_C1_H and Bin_OR = '0') then
         s_Energy_Bin_851 <= s_Energy_Bin_851 +'1';
		 Energy_Bin_Rdy_851 <= '1';
		else
		 s_Energy_Bin_851 <= s_Energy_Bin_851;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_851 <= '0';
      end if;
    end if;
  end process  Energy_Bin_851;   
  
  Energy_Bin_852 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_852   <=  (others =>'0');
	    Energy_Bin_Rdy_852 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E852_C1_L and PEAK_C1 <= s_E852_C1_H and Bin_OR = '0') then
         s_Energy_Bin_852 <= s_Energy_Bin_852 +'1';
		 Energy_Bin_Rdy_852 <= '1';
		else
		 s_Energy_Bin_852 <= s_Energy_Bin_852;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_852 <= '0';
      end if;
    end if;
  end process  Energy_Bin_852;   
  
  Energy_Bin_853 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_853   <=  (others =>'0');
	    Energy_Bin_Rdy_853 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E853_C1_L and PEAK_C1 <= s_E853_C1_H and Bin_OR = '0') then
         s_Energy_Bin_853 <= s_Energy_Bin_853 +'1';
		 Energy_Bin_Rdy_853 <= '1';
		else
		 s_Energy_Bin_853 <= s_Energy_Bin_853;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_853 <= '0';
      end if;
    end if;
  end process  Energy_Bin_853;   
  
  Energy_Bin_854 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_854   <=  (others =>'0');
		Energy_Bin_Rdy_854 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E854_C1_L and PEAK_C1 <= s_E854_C1_H and Bin_OR = '0') then
         s_Energy_Bin_854 <= s_Energy_Bin_854 +'1';
		 Energy_Bin_Rdy_854 <= '1';
		else
		 s_Energy_Bin_854 <= s_Energy_Bin_854;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_854 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_854;   
 
 
  Energy_Bin_855 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_855   <=  (others =>'0');
		Energy_Bin_Rdy_855 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E855_C1_L and PEAK_C1 <= s_E855_C1_H and Bin_OR = '0') then
         s_Energy_Bin_855 <= s_Energy_Bin_855 +'1';
		 Energy_Bin_Rdy_855 <= '1';
		else
		 s_Energy_Bin_855 <= s_Energy_Bin_855;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_855 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_855;  
 
  
  Energy_Bin_856 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_856   <=  (others =>'0');
		Energy_Bin_Rdy_856 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E856_C1_L and PEAK_C1 <= s_E856_C1_H and Bin_OR = '0') then
         s_Energy_Bin_856 <= s_Energy_Bin_856 +'1';
		 Energy_Bin_Rdy_856 <= '1';
		else
		 s_Energy_Bin_856 <= s_Energy_Bin_856;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_856 <= '0';
      end if;
    end if;
  end process  Energy_Bin_856;   
  
 Energy_Bin_857 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_857   <=  (others =>'0');
		Energy_Bin_Rdy_857 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E857_C1_L and PEAK_C1 <= s_E857_C1_H and Bin_OR = '0') then
         s_Energy_Bin_857 <= s_Energy_Bin_857 +'1';
		 Energy_Bin_Rdy_857 <= '1';
		else
		 s_Energy_Bin_857 <= s_Energy_Bin_857;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_857 <= '0';
      end if;
    end if;
  end process  Energy_Bin_857;   
  
  Energy_Bin_858 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_858   <=  (others =>'0');
		Energy_Bin_Rdy_858 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E858_C1_L and PEAK_C1 <= s_E858_C1_H and Bin_OR = '0') then
         s_Energy_Bin_858 <= s_Energy_Bin_858 +'1';
		 Energy_Bin_Rdy_858 <= '1';
		else
		 s_Energy_Bin_858 <= s_Energy_Bin_858;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_858 <= '0';
      end if;
    end if;
  end process  Energy_Bin_858;   
  
  Energy_Bin_859 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_859   <=  (others =>'0');
		Energy_Bin_Rdy_859 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E859_C1_L and PEAK_C1 <= s_E859_C1_H and Bin_OR = '0') then
         s_Energy_Bin_859 <= s_Energy_Bin_859 +'1';
		 Energy_Bin_Rdy_859 <= '1';
		else
		 s_Energy_Bin_859 <= s_Energy_Bin_859;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_859 <= '0';
      end if;
    end if;
  end process  Energy_Bin_859;           
  
     Energy_Bin_860 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_860   <=  (others =>'0');
		Energy_Bin_Rdy_860 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E860_C1_L and PEAK_C1 <= s_E860_C1_H and Bin_OR = '0') then
         s_Energy_Bin_860 <= s_Energy_Bin_860 +'1';
		 Energy_Bin_Rdy_860 <= '1';
		else
		 s_Energy_Bin_860 <= s_Energy_Bin_860;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_860 <= '0';
      end if;
    end if;
  end process  Energy_Bin_860;    
  
  Energy_Bin_861 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_861   <=  (others =>'0');
		Energy_Bin_Rdy_861 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E861_C1_L and PEAK_C1 <= s_E861_C1_H and Bin_OR = '0') then
         s_Energy_Bin_861 <= s_Energy_Bin_861 +'1';
		 Energy_Bin_Rdy_861 <= '1';
		else
		 s_Energy_Bin_861 <= s_Energy_Bin_861;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_861 <= '0';
      end if;
    end if;
  end process  Energy_Bin_861;   
  
  Energy_Bin_862 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_862   <=  (others =>'0');
	    Energy_Bin_Rdy_862 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E862_C1_L and PEAK_C1 <= s_E862_C1_H and Bin_OR = '0') then
         s_Energy_Bin_862 <= s_Energy_Bin_862 +'1';
		 Energy_Bin_Rdy_862 <= '1';
		else
		 s_Energy_Bin_862 <= s_Energy_Bin_862;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_862 <= '0';
      end if;
    end if;
  end process  Energy_Bin_862;   
  
  Energy_Bin_863 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_863   <=  (others =>'0');
	    Energy_Bin_Rdy_863 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E863_C1_L and PEAK_C1 <= s_E863_C1_H and Bin_OR = '0') then
         s_Energy_Bin_863 <= s_Energy_Bin_863 +'1';
		 Energy_Bin_Rdy_863 <= '1';
		else
		 s_Energy_Bin_863 <= s_Energy_Bin_863;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_863 <= '0';
      end if;
    end if;
  end process  Energy_Bin_863;   
  
  Energy_Bin_864 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_864   <=  (others =>'0');
		Energy_Bin_Rdy_864 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E864_C1_L and PEAK_C1 <= s_E864_C1_H and Bin_OR = '0') then
         s_Energy_Bin_864 <= s_Energy_Bin_864 +'1';
		 Energy_Bin_Rdy_864 <= '1';
		else
		 s_Energy_Bin_864 <= s_Energy_Bin_864;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_864 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_864;   
 
 
  Energy_Bin_865 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_865   <=  (others =>'0');
		Energy_Bin_Rdy_865 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E865_C1_L and PEAK_C1 <= s_E865_C1_H and Bin_OR = '0') then
         s_Energy_Bin_865 <= s_Energy_Bin_865 +'1';
		 Energy_Bin_Rdy_865 <= '1';
		else
		 s_Energy_Bin_865 <= s_Energy_Bin_865;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_865 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_865;  
 
  
  Energy_Bin_866 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_866   <=  (others =>'0');
		Energy_Bin_Rdy_866 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E866_C1_L and PEAK_C1 <= s_E866_C1_H and Bin_OR = '0') then
         s_Energy_Bin_866 <= s_Energy_Bin_866 +'1';
		 Energy_Bin_Rdy_866 <= '1';
		else
		 s_Energy_Bin_866 <= s_Energy_Bin_866;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_866 <= '0';
      end if;
    end if;
  end process  Energy_Bin_866;   
  
 Energy_Bin_867 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_867   <=  (others =>'0');
		Energy_Bin_Rdy_867 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E867_C1_L and PEAK_C1 <= s_E867_C1_H and Bin_OR = '0') then
         s_Energy_Bin_867 <= s_Energy_Bin_867 +'1';
		 Energy_Bin_Rdy_867 <= '1';
		else
		 s_Energy_Bin_867 <= s_Energy_Bin_867;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_867 <= '0';
      end if;
    end if;
  end process  Energy_Bin_867;   
  
  Energy_Bin_868 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_868   <=  (others =>'0');
		Energy_Bin_Rdy_868 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E868_C1_L and PEAK_C1 <= s_E868_C1_H and Bin_OR = '0') then
         s_Energy_Bin_868 <= s_Energy_Bin_868 +'1';
		 Energy_Bin_Rdy_868 <= '1';
		else
		 s_Energy_Bin_868 <= s_Energy_Bin_868;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_868 <= '0';
      end if;
    end if;
  end process  Energy_Bin_868;   
  
  Energy_Bin_869 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_869   <=  (others =>'0');
		Energy_Bin_Rdy_869 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E869_C1_L and PEAK_C1 <= s_E869_C1_H and Bin_OR = '0') then
         s_Energy_Bin_869 <= s_Energy_Bin_869 +'1';
		 Energy_Bin_Rdy_869 <= '1';
		else
		 s_Energy_Bin_869 <= s_Energy_Bin_869;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_869 <= '0';
      end if;
    end if;
  end process  Energy_Bin_869;         
  
     Energy_Bin_870 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_870   <=  (others =>'0');
		Energy_Bin_Rdy_870 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E870_C1_L and PEAK_C1 <= s_E870_C1_H and Bin_OR = '0') then
         s_Energy_Bin_870 <= s_Energy_Bin_870 +'1';
		 Energy_Bin_Rdy_870 <= '1';
		else
		 s_Energy_Bin_870 <= s_Energy_Bin_870;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_870 <= '0';
      end if;
    end if;
  end process  Energy_Bin_870;    
  
  Energy_Bin_871 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_871   <=  (others =>'0');
		Energy_Bin_Rdy_871 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E871_C1_L and PEAK_C1 <= s_E871_C1_H and Bin_OR = '0') then
         s_Energy_Bin_871 <= s_Energy_Bin_871 +'1';
		 Energy_Bin_Rdy_871 <= '1';
		else
		 s_Energy_Bin_871 <= s_Energy_Bin_871;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_871 <= '0';
      end if;
    end if;
  end process  Energy_Bin_871;   
  
  Energy_Bin_872 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_872   <=  (others =>'0');
	    Energy_Bin_Rdy_872 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E872_C1_L and PEAK_C1 <= s_E872_C1_H and Bin_OR = '0') then
         s_Energy_Bin_872 <= s_Energy_Bin_872 +'1';
		 Energy_Bin_Rdy_872 <= '1';
		else
		 s_Energy_Bin_872 <= s_Energy_Bin_872;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_872 <= '0';
      end if;
    end if;
  end process  Energy_Bin_872;   
  
  Energy_Bin_873 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_873   <=  (others =>'0');
	    Energy_Bin_Rdy_873 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E873_C1_L and PEAK_C1 <= s_E873_C1_H and Bin_OR = '0') then
         s_Energy_Bin_873 <= s_Energy_Bin_873 +'1';
		 Energy_Bin_Rdy_873 <= '1';
		else
		 s_Energy_Bin_873 <= s_Energy_Bin_873;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_873 <= '0';
      end if;
    end if;
  end process  Energy_Bin_873;   
  
  Energy_Bin_874 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_874   <=  (others =>'0');
		Energy_Bin_Rdy_874 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E874_C1_L and PEAK_C1 <= s_E874_C1_H and Bin_OR = '0') then
         s_Energy_Bin_874 <= s_Energy_Bin_874 +'1';
		 Energy_Bin_Rdy_874 <= '1';
		else
		 s_Energy_Bin_874 <= s_Energy_Bin_874;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_874 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_874;   
 
 
  Energy_Bin_875 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_875   <=  (others =>'0');
		Energy_Bin_Rdy_875 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E875_C1_L and PEAK_C1 <= s_E875_C1_H and Bin_OR = '0') then
         s_Energy_Bin_875 <= s_Energy_Bin_875 +'1';
		 Energy_Bin_Rdy_875 <= '1';
		else
		 s_Energy_Bin_875 <= s_Energy_Bin_875;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_875 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_875;  
 
  
  Energy_Bin_876 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_876   <=  (others =>'0');
		Energy_Bin_Rdy_876 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E876_C1_L and PEAK_C1 <= s_E876_C1_H and Bin_OR = '0') then
         s_Energy_Bin_876 <= s_Energy_Bin_876 +'1';
		 Energy_Bin_Rdy_876 <= '1';
		else
		 s_Energy_Bin_876 <= s_Energy_Bin_876;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_876 <= '0';
      end if;
    end if;
  end process  Energy_Bin_876;   
  
 Energy_Bin_877 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_877   <=  (others =>'0');
		Energy_Bin_Rdy_877 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E877_C1_L and PEAK_C1 <= s_E877_C1_H and Bin_OR = '0') then
         s_Energy_Bin_877 <= s_Energy_Bin_877 +'1';
		 Energy_Bin_Rdy_877 <= '1';
		else
		 s_Energy_Bin_877 <= s_Energy_Bin_877;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_877 <= '0';
      end if;
    end if;
  end process  Energy_Bin_877;   
  
  Energy_Bin_878 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_878   <=  (others =>'0');
		Energy_Bin_Rdy_878 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E878_C1_L and PEAK_C1 <= s_E878_C1_H and Bin_OR = '0') then
         s_Energy_Bin_878 <= s_Energy_Bin_878 +'1';
		 Energy_Bin_Rdy_878 <= '1';
		else
		 s_Energy_Bin_878 <= s_Energy_Bin_878;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_878 <= '0';
      end if;
    end if;
  end process  Energy_Bin_878;   
  
  Energy_Bin_879 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_879   <=  (others =>'0');
		Energy_Bin_Rdy_879 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E879_C1_L and PEAK_C1 <= s_E879_C1_H and Bin_OR = '0') then
         s_Energy_Bin_879 <= s_Energy_Bin_879 +'1';
		 Energy_Bin_Rdy_879 <= '1';
		else
		 s_Energy_Bin_879 <= s_Energy_Bin_879;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_879 <= '0';
      end if;
    end if;
  end process  Energy_Bin_879;       
  
     Energy_Bin_880 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_880   <=  (others =>'0');
		Energy_Bin_Rdy_880 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E880_C1_L and PEAK_C1 <= s_E880_C1_H and Bin_OR = '0') then
         s_Energy_Bin_880 <= s_Energy_Bin_880 +'1';
		 Energy_Bin_Rdy_880 <= '1';
		else
		 s_Energy_Bin_880 <= s_Energy_Bin_880;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_880 <= '0';
      end if;
    end if;
  end process  Energy_Bin_880;    
  
  Energy_Bin_881 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_881   <=  (others =>'0');
		Energy_Bin_Rdy_881 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E881_C1_L and PEAK_C1 <= s_E881_C1_H and Bin_OR = '0') then
         s_Energy_Bin_881 <= s_Energy_Bin_881 +'1';
		 Energy_Bin_Rdy_881 <= '1';
		else
		 s_Energy_Bin_881 <= s_Energy_Bin_881;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_881 <= '0';
      end if;
    end if;
  end process  Energy_Bin_881;   
  
  Energy_Bin_882 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_882   <=  (others =>'0');
	    Energy_Bin_Rdy_882 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E882_C1_L and PEAK_C1 <= s_E882_C1_H and Bin_OR = '0') then
         s_Energy_Bin_882 <= s_Energy_Bin_882 +'1';
		 Energy_Bin_Rdy_882 <= '1';
		else
		 s_Energy_Bin_882 <= s_Energy_Bin_882;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_882 <= '0';
      end if;
    end if;
  end process  Energy_Bin_882;   
  
  Energy_Bin_883 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_883   <=  (others =>'0');
	    Energy_Bin_Rdy_883 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E883_C1_L and PEAK_C1 <= s_E883_C1_H and Bin_OR = '0') then
         s_Energy_Bin_883 <= s_Energy_Bin_883 +'1';
		 Energy_Bin_Rdy_883 <= '1';
		else
		 s_Energy_Bin_883 <= s_Energy_Bin_883;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_883 <= '0';
      end if;
    end if;
  end process  Energy_Bin_883;   
  
  Energy_Bin_884 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_884   <=  (others =>'0');
		Energy_Bin_Rdy_884 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E884_C1_L and PEAK_C1 <= s_E884_C1_H and Bin_OR = '0') then
         s_Energy_Bin_884 <= s_Energy_Bin_884 +'1';
		 Energy_Bin_Rdy_884 <= '1';
		else
		 s_Energy_Bin_884 <= s_Energy_Bin_884;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_884 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_884;   
 
 
  Energy_Bin_885 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_885   <=  (others =>'0');
		Energy_Bin_Rdy_885 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E885_C1_L and PEAK_C1 <= s_E885_C1_H and Bin_OR = '0') then
         s_Energy_Bin_885 <= s_Energy_Bin_885 +'1';
		 Energy_Bin_Rdy_885 <= '1';
		else
		 s_Energy_Bin_885 <= s_Energy_Bin_885;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_885 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_885;  
 
  
  Energy_Bin_886 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_886   <=  (others =>'0');
		Energy_Bin_Rdy_886 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E886_C1_L and PEAK_C1 <= s_E886_C1_H and Bin_OR = '0') then
         s_Energy_Bin_886 <= s_Energy_Bin_886 +'1';
		 Energy_Bin_Rdy_886 <= '1';
		else
		 s_Energy_Bin_886 <= s_Energy_Bin_886;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_886 <= '0';
      end if;
    end if;
  end process  Energy_Bin_886;   
  
 Energy_Bin_887 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_887   <=  (others =>'0');
		Energy_Bin_Rdy_887 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E887_C1_L and PEAK_C1 <= s_E887_C1_H and Bin_OR = '0') then
         s_Energy_Bin_887 <= s_Energy_Bin_887 +'1';
		 Energy_Bin_Rdy_887 <= '1';
		else
		 s_Energy_Bin_887 <= s_Energy_Bin_887;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_887 <= '0';
      end if;
    end if;
  end process  Energy_Bin_887;   
  
  Energy_Bin_888 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_888   <=  (others =>'0');
		Energy_Bin_Rdy_888 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E888_C1_L and PEAK_C1 <= s_E888_C1_H and Bin_OR = '0') then
         s_Energy_Bin_888 <= s_Energy_Bin_888 +'1';
		 Energy_Bin_Rdy_888 <= '1';
		else
		 s_Energy_Bin_888 <= s_Energy_Bin_888;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_888 <= '0';
      end if;
    end if;
  end process  Energy_Bin_888;   
  
  Energy_Bin_889 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_889   <=  (others =>'0');
		Energy_Bin_Rdy_889 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E889_C1_L and PEAK_C1 <= s_E889_C1_H and Bin_OR = '0') then
         s_Energy_Bin_889 <= s_Energy_Bin_889 +'1';
		 Energy_Bin_Rdy_889 <= '1';
		else
		 s_Energy_Bin_889 <= s_Energy_Bin_889;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_889 <= '0';
      end if;
    end if;
  end process  Energy_Bin_889;      
  
     Energy_Bin_890 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_890   <=  (others =>'0');
		Energy_Bin_Rdy_890 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E890_C1_L and PEAK_C1 <= s_E890_C1_H and Bin_OR = '0') then
         s_Energy_Bin_890 <= s_Energy_Bin_890 +'1';
		 Energy_Bin_Rdy_890 <= '1';
		else
		 s_Energy_Bin_890 <= s_Energy_Bin_890;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_890 <= '0';
      end if;
    end if;
  end process  Energy_Bin_890;    
  
  Energy_Bin_891 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_891   <=  (others =>'0');
		Energy_Bin_Rdy_891 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E891_C1_L and PEAK_C1 <= s_E891_C1_H and Bin_OR = '0') then
         s_Energy_Bin_891 <= s_Energy_Bin_891 +'1';
		 Energy_Bin_Rdy_891 <= '1';
		else
		 s_Energy_Bin_891 <= s_Energy_Bin_891;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_891 <= '0';
      end if;
    end if;
  end process  Energy_Bin_891;   
  
  Energy_Bin_892 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_892   <=  (others =>'0');
	    Energy_Bin_Rdy_892 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E892_C1_L and PEAK_C1 <= s_E892_C1_H and Bin_OR = '0') then
         s_Energy_Bin_892 <= s_Energy_Bin_892 +'1';
		 Energy_Bin_Rdy_892 <= '1';
		else
		 s_Energy_Bin_892 <= s_Energy_Bin_892;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_892 <= '0';
      end if;
    end if;
  end process  Energy_Bin_892;   
  
  Energy_Bin_893 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_893   <=  (others =>'0');
	    Energy_Bin_Rdy_893 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E893_C1_L and PEAK_C1 <= s_E893_C1_H and Bin_OR = '0') then
         s_Energy_Bin_893 <= s_Energy_Bin_893 +'1';
		 Energy_Bin_Rdy_893 <= '1';
		else
		 s_Energy_Bin_893 <= s_Energy_Bin_893;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_893 <= '0';
      end if;
    end if;
  end process  Energy_Bin_893;   
  
  Energy_Bin_894 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_894   <=  (others =>'0');
		Energy_Bin_Rdy_894 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E894_C1_L and PEAK_C1 <= s_E894_C1_H and Bin_OR = '0') then
         s_Energy_Bin_894 <= s_Energy_Bin_894 +'1';
		 Energy_Bin_Rdy_894 <= '1';
		else
		 s_Energy_Bin_894 <= s_Energy_Bin_894;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_894 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_894;   
 
 
  Energy_Bin_895 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_895   <=  (others =>'0');
		Energy_Bin_Rdy_895 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E895_C1_L and PEAK_C1 <= s_E895_C1_H and Bin_OR = '0') then
         s_Energy_Bin_895 <= s_Energy_Bin_895 +'1';
		 Energy_Bin_Rdy_895 <= '1';
		else
		 s_Energy_Bin_895 <= s_Energy_Bin_895;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_895 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_895;  
 
  
  Energy_Bin_896 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_896   <=  (others =>'0');
		Energy_Bin_Rdy_896 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E896_C1_L and PEAK_C1 <= s_E896_C1_H and Bin_OR = '0') then
         s_Energy_Bin_896 <= s_Energy_Bin_896 +'1';
		 Energy_Bin_Rdy_896 <= '1';
		else
		 s_Energy_Bin_896 <= s_Energy_Bin_896;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_896 <= '0';
      end if;
    end if;
  end process  Energy_Bin_896;   
  
 Energy_Bin_897 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_897   <=  (others =>'0');
		Energy_Bin_Rdy_897 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E897_C1_L and PEAK_C1 <= s_E897_C1_H and Bin_OR = '0') then
         s_Energy_Bin_897 <= s_Energy_Bin_897 +'1';
		 Energy_Bin_Rdy_897 <= '1';
		else
		 s_Energy_Bin_897 <= s_Energy_Bin_897;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_897 <= '0';
      end if;
    end if;
  end process  Energy_Bin_897;   
  
  Energy_Bin_898 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_898   <=  (others =>'0');
		Energy_Bin_Rdy_898 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E898_C1_L and PEAK_C1 <= s_E898_C1_H and Bin_OR = '0') then
         s_Energy_Bin_898 <= s_Energy_Bin_898 +'1';
		 Energy_Bin_Rdy_898 <= '1';
		else
		 s_Energy_Bin_898 <= s_Energy_Bin_898;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_898 <= '0';
      end if;
    end if;
  end process  Energy_Bin_898;   
  
  Energy_Bin_899 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_899   <=  (others =>'0');
		Energy_Bin_Rdy_899 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E899_C1_L and PEAK_C1 <= s_E899_C1_H and Bin_OR = '0') then
         s_Energy_Bin_899 <= s_Energy_Bin_899 +'1';
		 Energy_Bin_Rdy_899 <= '1';
		else
		 s_Energy_Bin_899 <= s_Energy_Bin_899;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_899 <= '0';
      end if;
    end if;
  end process  Energy_Bin_899;   

    Energy_Bin_900 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_900   <=  (others =>'0');
		Energy_Bin_Rdy_900 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E900_C1_L and PEAK_C1 <= s_E900_C1_H and Bin_OR = '0') then
         s_Energy_Bin_900 <= s_Energy_Bin_900 +'1';
		 Energy_Bin_Rdy_900 <= '1';
		else
		 s_Energy_Bin_900 <= s_Energy_Bin_900;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_900 <= '0';
      end if;
    end if;
  end process  Energy_Bin_900;    
  
  Energy_Bin_901 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_901   <=  (others =>'0');
		Energy_Bin_Rdy_901 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E901_C1_L and PEAK_C1 <= s_E901_C1_H and Bin_OR = '0') then
         s_Energy_Bin_901 <= s_Energy_Bin_901 +'1';
		 Energy_Bin_Rdy_901 <= '1';
		else
		 s_Energy_Bin_901 <= s_Energy_Bin_901;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_901 <= '0';
      end if;
    end if;
  end process  Energy_Bin_901;   
  
  Energy_Bin_902 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_902   <=  (others =>'0');
	    Energy_Bin_Rdy_902 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E902_C1_L and PEAK_C1 <= s_E902_C1_H and Bin_OR = '0') then
         s_Energy_Bin_902 <= s_Energy_Bin_902 +'1';
		 Energy_Bin_Rdy_902 <= '1';
		else
		 s_Energy_Bin_902 <= s_Energy_Bin_902;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_902 <= '0';
      end if;
    end if;
  end process  Energy_Bin_902;   
  
  Energy_Bin_903 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_903   <=  (others =>'0');
	    Energy_Bin_Rdy_903 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E903_C1_L and PEAK_C1 <= s_E903_C1_H and Bin_OR = '0') then
         s_Energy_Bin_903 <= s_Energy_Bin_903 +'1';
		 Energy_Bin_Rdy_903 <= '1';
		else
		 s_Energy_Bin_903 <= s_Energy_Bin_903;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_903 <= '0';
      end if;
    end if;
  end process  Energy_Bin_903;   
  
  Energy_Bin_904 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_904   <=  (others =>'0');
		Energy_Bin_Rdy_904 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E904_C1_L and PEAK_C1 <= s_E904_C1_H and Bin_OR = '0') then
         s_Energy_Bin_904 <= s_Energy_Bin_904 +'1';
		 Energy_Bin_Rdy_904 <= '1';
		else
		 s_Energy_Bin_904 <= s_Energy_Bin_904;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_904 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_904;   
 
 
  Energy_Bin_905 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_905   <=  (others =>'0');
		Energy_Bin_Rdy_905 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E905_C1_L and PEAK_C1 <= s_E905_C1_H and Bin_OR = '0') then
         s_Energy_Bin_905 <= s_Energy_Bin_905 +'1';
		 Energy_Bin_Rdy_905 <= '1';
		else
		 s_Energy_Bin_905 <= s_Energy_Bin_905;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_905 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_905;  
 
  
  Energy_Bin_906 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_906   <=  (others =>'0');
		Energy_Bin_Rdy_906 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E906_C1_L and PEAK_C1 <= s_E906_C1_H and Bin_OR = '0') then
         s_Energy_Bin_906 <= s_Energy_Bin_906 +'1';
		 Energy_Bin_Rdy_906 <= '1';
		else
		 s_Energy_Bin_906 <= s_Energy_Bin_906;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_906 <= '0';
      end if;
    end if;
  end process  Energy_Bin_906;   
  
 Energy_Bin_907 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_907   <=  (others =>'0');
		Energy_Bin_Rdy_907 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E907_C1_L and PEAK_C1 <= s_E907_C1_H and Bin_OR = '0') then
         s_Energy_Bin_907 <= s_Energy_Bin_907 +'1';
		 Energy_Bin_Rdy_907 <= '1';
		else
		 s_Energy_Bin_907 <= s_Energy_Bin_907;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_907 <= '0';
      end if;
    end if;
  end process  Energy_Bin_907;   
  
  Energy_Bin_908 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_908   <=  (others =>'0');
		Energy_Bin_Rdy_908 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E908_C1_L and PEAK_C1 <= s_E908_C1_H and Bin_OR = '0') then
         s_Energy_Bin_908 <= s_Energy_Bin_908 +'1';
		 Energy_Bin_Rdy_908 <= '1';
		else
		 s_Energy_Bin_908 <= s_Energy_Bin_908;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_908 <= '0';
      end if;
    end if;
  end process  Energy_Bin_908;   
  
  Energy_Bin_909 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_909   <=  (others =>'0');
		Energy_Bin_Rdy_909 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E909_C1_L and PEAK_C1 <= s_E909_C1_H and Bin_OR = '0') then
         s_Energy_Bin_909 <= s_Energy_Bin_909 +'1';
		 Energy_Bin_Rdy_909 <= '1';
		else
		 s_Energy_Bin_909 <= s_Energy_Bin_909;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_909 <= '0';
      end if;
    end if;
  end process  Energy_Bin_909;      
  
     Energy_Bin_910 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_910   <=  (others =>'0');
		Energy_Bin_Rdy_910 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E910_C1_L and PEAK_C1 <= s_E910_C1_H and Bin_OR = '0') then
         s_Energy_Bin_910 <= s_Energy_Bin_910 +'1';
		 Energy_Bin_Rdy_910 <= '1';
		else
		 s_Energy_Bin_910 <= s_Energy_Bin_910;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_910 <= '0';
      end if;
    end if;
  end process  Energy_Bin_910;    
  
  Energy_Bin_911 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_911   <=  (others =>'0');
		Energy_Bin_Rdy_911 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E911_C1_L and PEAK_C1 <= s_E911_C1_H and Bin_OR = '0') then
         s_Energy_Bin_911 <= s_Energy_Bin_911 +'1';
		 Energy_Bin_Rdy_911 <= '1';
		else
		 s_Energy_Bin_911 <= s_Energy_Bin_911;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_911 <= '0';
      end if;
    end if;
  end process  Energy_Bin_911;   
  
  Energy_Bin_912 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_912   <=  (others =>'0');
	    Energy_Bin_Rdy_912 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E912_C1_L and PEAK_C1 <= s_E912_C1_H and Bin_OR = '0') then
         s_Energy_Bin_912 <= s_Energy_Bin_912 +'1';
		 Energy_Bin_Rdy_912 <= '1';
		else
		 s_Energy_Bin_912 <= s_Energy_Bin_912;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_912 <= '0';
      end if;
    end if;
  end process  Energy_Bin_912;   
  
  Energy_Bin_913 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_913   <=  (others =>'0');
	    Energy_Bin_Rdy_913 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E913_C1_L and PEAK_C1 <= s_E913_C1_H and Bin_OR = '0') then
         s_Energy_Bin_913 <= s_Energy_Bin_913 +'1';
		 Energy_Bin_Rdy_913 <= '1';
		else
		 s_Energy_Bin_913 <= s_Energy_Bin_913;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_913 <= '0';
      end if;
    end if;
  end process  Energy_Bin_913;   
  
  Energy_Bin_914 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_914   <=  (others =>'0');
		Energy_Bin_Rdy_914 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E914_C1_L and PEAK_C1 <= s_E914_C1_H and Bin_OR = '0') then
         s_Energy_Bin_914 <= s_Energy_Bin_914 +'1';
		 Energy_Bin_Rdy_914 <= '1';
		else
		 s_Energy_Bin_914 <= s_Energy_Bin_914;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_914 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_914;   
 
 
  Energy_Bin_915 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_915   <=  (others =>'0');
		Energy_Bin_Rdy_915 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E915_C1_L and PEAK_C1 <= s_E915_C1_H and Bin_OR = '0') then
         s_Energy_Bin_915 <= s_Energy_Bin_915 +'1';
		 Energy_Bin_Rdy_915 <= '1';
		else
		 s_Energy_Bin_915 <= s_Energy_Bin_915;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_915 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_915;  
 
  
  Energy_Bin_916 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_916   <=  (others =>'0');
		Energy_Bin_Rdy_916 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E916_C1_L and PEAK_C1 <= s_E916_C1_H and Bin_OR = '0') then
         s_Energy_Bin_916 <= s_Energy_Bin_916 +'1';
		 Energy_Bin_Rdy_916 <= '1';
		else
		 s_Energy_Bin_916 <= s_Energy_Bin_916;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_916 <= '0';
      end if;
    end if;
  end process  Energy_Bin_916;   
  
 Energy_Bin_917 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_917   <=  (others =>'0');
		Energy_Bin_Rdy_917 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E917_C1_L and PEAK_C1 <= s_E917_C1_H and Bin_OR = '0') then
         s_Energy_Bin_917 <= s_Energy_Bin_917 +'1';
		 Energy_Bin_Rdy_917 <= '1';
		else
		 s_Energy_Bin_917 <= s_Energy_Bin_917;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_917 <= '0';
      end if;
    end if;
  end process  Energy_Bin_917;   
  
  Energy_Bin_918 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_918   <=  (others =>'0');
		Energy_Bin_Rdy_918 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E918_C1_L and PEAK_C1 <= s_E918_C1_H and Bin_OR = '0') then
         s_Energy_Bin_918 <= s_Energy_Bin_918 +'1';
		 Energy_Bin_Rdy_918 <= '1';
		else
		 s_Energy_Bin_918 <= s_Energy_Bin_918;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_918 <= '0';
      end if;
    end if;
  end process  Energy_Bin_918;   
  
  Energy_Bin_919 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_919   <=  (others =>'0');
		Energy_Bin_Rdy_919 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E919_C1_L and PEAK_C1 <= s_E919_C1_H and Bin_OR = '0') then
         s_Energy_Bin_919 <= s_Energy_Bin_919 +'1';
		 Energy_Bin_Rdy_919 <= '1';
		else
		 s_Energy_Bin_919 <= s_Energy_Bin_919;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_919 <= '0';
      end if;
    end if;
  end process  Energy_Bin_919;       
  
     Energy_Bin_920 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_920   <=  (others =>'0');
		Energy_Bin_Rdy_920 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E920_C1_L and PEAK_C1 <= s_E920_C1_H and Bin_OR = '0') then
         s_Energy_Bin_920 <= s_Energy_Bin_920 +'1';
		 Energy_Bin_Rdy_920 <= '1';
		else
		 s_Energy_Bin_920 <= s_Energy_Bin_920;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_920 <= '0';
      end if;
    end if;
  end process  Energy_Bin_920;    
  
  Energy_Bin_921 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_921   <=  (others =>'0');
		Energy_Bin_Rdy_921 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E921_C1_L and PEAK_C1 <= s_E921_C1_H and Bin_OR = '0') then
         s_Energy_Bin_921 <= s_Energy_Bin_921 +'1';
		 Energy_Bin_Rdy_921 <= '1';
		else
		 s_Energy_Bin_921 <= s_Energy_Bin_921;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_921 <= '0';
      end if;
    end if;
  end process  Energy_Bin_921;   
  
  Energy_Bin_922 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_922   <=  (others =>'0');
	    Energy_Bin_Rdy_922 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E922_C1_L and PEAK_C1 <= s_E922_C1_H and Bin_OR = '0') then
         s_Energy_Bin_922 <= s_Energy_Bin_922 +'1';
		 Energy_Bin_Rdy_922 <= '1';
		else
		 s_Energy_Bin_922 <= s_Energy_Bin_922;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_922 <= '0';
      end if;
    end if;
  end process  Energy_Bin_922;   
  
  Energy_Bin_923 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_923   <=  (others =>'0');
	    Energy_Bin_Rdy_923 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E923_C1_L and PEAK_C1 <= s_E923_C1_H and Bin_OR = '0') then
         s_Energy_Bin_923 <= s_Energy_Bin_923 +'1';
		 Energy_Bin_Rdy_923 <= '1';
		else
		 s_Energy_Bin_923 <= s_Energy_Bin_923;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_923 <= '0';
      end if;
    end if;
  end process  Energy_Bin_923;   
  
  Energy_Bin_924 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_924   <=  (others =>'0');
		Energy_Bin_Rdy_924 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E924_C1_L and PEAK_C1 <= s_E924_C1_H and Bin_OR = '0') then
         s_Energy_Bin_924 <= s_Energy_Bin_924 +'1';
		 Energy_Bin_Rdy_924 <= '1';
		else
		 s_Energy_Bin_924 <= s_Energy_Bin_924;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_924 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_924;   
 
 
  Energy_Bin_925 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_925   <=  (others =>'0');
		Energy_Bin_Rdy_925 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E925_C1_L and PEAK_C1 <= s_E925_C1_H and Bin_OR = '0') then
         s_Energy_Bin_925 <= s_Energy_Bin_925 +'1';
		 Energy_Bin_Rdy_925 <= '1';
		else
		 s_Energy_Bin_925 <= s_Energy_Bin_925;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_925 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_925;  
 
  
  Energy_Bin_926 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_926   <=  (others =>'0');
		Energy_Bin_Rdy_926 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E926_C1_L and PEAK_C1 <= s_E926_C1_H and Bin_OR = '0') then
         s_Energy_Bin_926 <= s_Energy_Bin_926 +'1';
		 Energy_Bin_Rdy_926 <= '1';
		else
		 s_Energy_Bin_926 <= s_Energy_Bin_926;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_926 <= '0';
      end if;
    end if;
  end process  Energy_Bin_926;   
  
 Energy_Bin_927 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_927   <=  (others =>'0');
		Energy_Bin_Rdy_927 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E927_C1_L and PEAK_C1 <= s_E927_C1_H and Bin_OR = '0') then
         s_Energy_Bin_927 <= s_Energy_Bin_927 +'1';
		 Energy_Bin_Rdy_927 <= '1';
		else
		 s_Energy_Bin_927 <= s_Energy_Bin_927;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_927 <= '0';
      end if;
    end if;
  end process  Energy_Bin_927;   
  
  Energy_Bin_928 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_928   <=  (others =>'0');
		Energy_Bin_Rdy_928 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E928_C1_L and PEAK_C1 <= s_E928_C1_H and Bin_OR = '0') then
         s_Energy_Bin_928 <= s_Energy_Bin_928 +'1';
		 Energy_Bin_Rdy_928 <= '1';
		else
		 s_Energy_Bin_928 <= s_Energy_Bin_928;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_928 <= '0';
      end if;
    end if;
  end process  Energy_Bin_928;   
  
  Energy_Bin_929 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_929   <=  (others =>'0');
		Energy_Bin_Rdy_929 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E929_C1_L and PEAK_C1 <= s_E929_C1_H and Bin_OR = '0') then
         s_Energy_Bin_929 <= s_Energy_Bin_929 +'1';
		 Energy_Bin_Rdy_929 <= '1';
		else
		 s_Energy_Bin_929 <= s_Energy_Bin_929;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_929 <= '0';
      end if;
    end if;
  end process  Energy_Bin_929;        
  
     Energy_Bin_930 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_930   <=  (others =>'0');
		Energy_Bin_Rdy_930 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E930_C1_L and PEAK_C1 <= s_E930_C1_H and Bin_OR = '0') then
         s_Energy_Bin_930 <= s_Energy_Bin_930 +'1';
		 Energy_Bin_Rdy_930 <= '1';
		else
		 s_Energy_Bin_930 <= s_Energy_Bin_930;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_930 <= '0';
      end if;
    end if;
  end process  Energy_Bin_930;    
  
  Energy_Bin_931 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_931   <=  (others =>'0');
		Energy_Bin_Rdy_931 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E931_C1_L and PEAK_C1 <= s_E931_C1_H and Bin_OR = '0') then
         s_Energy_Bin_931 <= s_Energy_Bin_931 +'1';
		 Energy_Bin_Rdy_931 <= '1';
		else
		 s_Energy_Bin_931 <= s_Energy_Bin_931;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_931 <= '0';
      end if;
    end if;
  end process  Energy_Bin_931;   
  
  Energy_Bin_932 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_932   <=  (others =>'0');
	    Energy_Bin_Rdy_932 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E932_C1_L and PEAK_C1 <= s_E932_C1_H and Bin_OR = '0') then
         s_Energy_Bin_932 <= s_Energy_Bin_932 +'1';
		 Energy_Bin_Rdy_932 <= '1';
		else
		 s_Energy_Bin_932 <= s_Energy_Bin_932;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_932 <= '0';
      end if;
    end if;
  end process  Energy_Bin_932;   
  
  Energy_Bin_933 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_933   <=  (others =>'0');
	    Energy_Bin_Rdy_933 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E933_C1_L and PEAK_C1 <= s_E933_C1_H and Bin_OR = '0') then
         s_Energy_Bin_933 <= s_Energy_Bin_933 +'1';
		 Energy_Bin_Rdy_933 <= '1';
		else
		 s_Energy_Bin_933 <= s_Energy_Bin_933;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_933 <= '0';
      end if;
    end if;
  end process  Energy_Bin_933;   
  
  Energy_Bin_934 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_934   <=  (others =>'0');
		Energy_Bin_Rdy_934 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E934_C1_L and PEAK_C1 <= s_E934_C1_H and Bin_OR = '0') then
         s_Energy_Bin_934 <= s_Energy_Bin_934 +'1';
		 Energy_Bin_Rdy_934 <= '1';
		else
		 s_Energy_Bin_934 <= s_Energy_Bin_934;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_934 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_934;   
 
 
  Energy_Bin_935 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_935   <=  (others =>'0');
		Energy_Bin_Rdy_935 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E935_C1_L and PEAK_C1 <= s_E935_C1_H and Bin_OR = '0') then
         s_Energy_Bin_935 <= s_Energy_Bin_935 +'1';
		 Energy_Bin_Rdy_935 <= '1';
		else
		 s_Energy_Bin_935 <= s_Energy_Bin_935;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_935 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_935;  
 
  
  Energy_Bin_936 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_936   <=  (others =>'0');
		Energy_Bin_Rdy_936 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E936_C1_L and PEAK_C1 <= s_E936_C1_H and Bin_OR = '0') then
         s_Energy_Bin_936 <= s_Energy_Bin_936 +'1';
		 Energy_Bin_Rdy_936 <= '1';
		else
		 s_Energy_Bin_936 <= s_Energy_Bin_936;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_936 <= '0';
      end if;
    end if;
  end process  Energy_Bin_936;   
  
 Energy_Bin_937 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_937   <=  (others =>'0');
		Energy_Bin_Rdy_937 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E937_C1_L and PEAK_C1 <= s_E937_C1_H and Bin_OR = '0') then
         s_Energy_Bin_937 <= s_Energy_Bin_937 +'1';
		 Energy_Bin_Rdy_937 <= '1';
		else
		 s_Energy_Bin_937 <= s_Energy_Bin_937;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_937 <= '0';
      end if;
    end if;
  end process  Energy_Bin_937;   
  
  Energy_Bin_938 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_938   <=  (others =>'0');
		Energy_Bin_Rdy_938 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E938_C1_L and PEAK_C1 <= s_E938_C1_H and Bin_OR = '0') then
         s_Energy_Bin_938 <= s_Energy_Bin_938 +'1';
		 Energy_Bin_Rdy_938 <= '1';
		else
		 s_Energy_Bin_938 <= s_Energy_Bin_938;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_938 <= '0';
      end if;
    end if;
  end process  Energy_Bin_938;   
  
  Energy_Bin_939 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_939   <=  (others =>'0');
		Energy_Bin_Rdy_939 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E939_C1_L and PEAK_C1 <= s_E939_C1_H and Bin_OR = '0') then
         s_Energy_Bin_939 <= s_Energy_Bin_939 +'1';
		 Energy_Bin_Rdy_939 <= '1';
		else
		 s_Energy_Bin_939 <= s_Energy_Bin_939;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_939 <= '0';
      end if;
    end if;
  end process  Energy_Bin_939;         
  
     Energy_Bin_940 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_940   <=  (others =>'0');
		Energy_Bin_Rdy_940 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E940_C1_L and PEAK_C1 <= s_E940_C1_H and Bin_OR = '0') then
         s_Energy_Bin_940 <= s_Energy_Bin_940 +'1';
		 Energy_Bin_Rdy_940 <= '1';
		else
		 s_Energy_Bin_940 <= s_Energy_Bin_940;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_940 <= '0';
      end if;
    end if;
  end process  Energy_Bin_940;    
  
  Energy_Bin_941 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_941   <=  (others =>'0');
		Energy_Bin_Rdy_941 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E941_C1_L and PEAK_C1 <= s_E941_C1_H and Bin_OR = '0') then
         s_Energy_Bin_941 <= s_Energy_Bin_941 +'1';
		 Energy_Bin_Rdy_941 <= '1';
		else
		 s_Energy_Bin_941 <= s_Energy_Bin_941;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_941 <= '0';
      end if;
    end if;
  end process  Energy_Bin_941;   
  
  Energy_Bin_942 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_942   <=  (others =>'0');
	    Energy_Bin_Rdy_942 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E942_C1_L and PEAK_C1 <= s_E942_C1_H and Bin_OR = '0') then
         s_Energy_Bin_942 <= s_Energy_Bin_942 +'1';
		 Energy_Bin_Rdy_942 <= '1';
		else
		 s_Energy_Bin_942 <= s_Energy_Bin_942;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_942 <= '0';
      end if;
    end if;
  end process  Energy_Bin_942;   
  
  Energy_Bin_943 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_943   <=  (others =>'0');
	    Energy_Bin_Rdy_943 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E943_C1_L and PEAK_C1 <= s_E943_C1_H and Bin_OR = '0') then
         s_Energy_Bin_943 <= s_Energy_Bin_943 +'1';
		 Energy_Bin_Rdy_943 <= '1';
		else
		 s_Energy_Bin_943 <= s_Energy_Bin_943;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_943 <= '0';
      end if;
    end if;
  end process  Energy_Bin_943;   
  
  Energy_Bin_944 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_944   <=  (others =>'0');
		Energy_Bin_Rdy_944 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E944_C1_L and PEAK_C1 <= s_E944_C1_H and Bin_OR = '0') then
         s_Energy_Bin_944 <= s_Energy_Bin_944 +'1';
		 Energy_Bin_Rdy_944 <= '1';
		else
		 s_Energy_Bin_944 <= s_Energy_Bin_944;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_944 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_944;   
 
 
  Energy_Bin_945 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_945   <=  (others =>'0');
		Energy_Bin_Rdy_945 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E945_C1_L and PEAK_C1 <= s_E945_C1_H and Bin_OR = '0') then
         s_Energy_Bin_945 <= s_Energy_Bin_945 +'1';
		 Energy_Bin_Rdy_945 <= '1';
		else
		 s_Energy_Bin_945 <= s_Energy_Bin_945;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_945 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_945;  
 
  
  Energy_Bin_946 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_946   <=  (others =>'0');
		Energy_Bin_Rdy_946 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E946_C1_L and PEAK_C1 <= s_E946_C1_H and Bin_OR = '0') then
         s_Energy_Bin_946 <= s_Energy_Bin_946 +'1';
		 Energy_Bin_Rdy_946 <= '1';
		else
		 s_Energy_Bin_946 <= s_Energy_Bin_946;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_946 <= '0';
      end if;
    end if;
  end process  Energy_Bin_946;   
  
 Energy_Bin_947 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_947   <=  (others =>'0');
		Energy_Bin_Rdy_947 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E947_C1_L and PEAK_C1 <= s_E947_C1_H and Bin_OR = '0') then
         s_Energy_Bin_947 <= s_Energy_Bin_947 +'1';
		 Energy_Bin_Rdy_947 <= '1';
		else
		 s_Energy_Bin_947 <= s_Energy_Bin_947;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_947 <= '0';
      end if;
    end if;
  end process  Energy_Bin_947;   
  
  Energy_Bin_948 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_948   <=  (others =>'0');
		Energy_Bin_Rdy_948 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E948_C1_L and PEAK_C1 <= s_E948_C1_H and Bin_OR = '0') then
         s_Energy_Bin_948 <= s_Energy_Bin_948 +'1';
		 Energy_Bin_Rdy_948 <= '1';
		else
		 s_Energy_Bin_948 <= s_Energy_Bin_948;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_948 <= '0';
      end if;
    end if;
  end process  Energy_Bin_948;   
  
  Energy_Bin_949 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_949   <=  (others =>'0');
		Energy_Bin_Rdy_949 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E949_C1_L and PEAK_C1 <= s_E949_C1_H and Bin_OR = '0') then
         s_Energy_Bin_949 <= s_Energy_Bin_949 +'1';
		 Energy_Bin_Rdy_949 <= '1';
		else
		 s_Energy_Bin_949 <= s_Energy_Bin_949;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_949 <= '0';
      end if;
    end if;
  end process  Energy_Bin_949;          
  
  
     Energy_Bin_950 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_950   <=  (others =>'0');
		Energy_Bin_Rdy_950 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E950_C1_L and PEAK_C1 <= s_E950_C1_H and Bin_OR = '0') then
         s_Energy_Bin_950 <= s_Energy_Bin_950 +'1';
		 Energy_Bin_Rdy_950 <= '1';
		else
		 s_Energy_Bin_950 <= s_Energy_Bin_950;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_950 <= '0';
      end if;
    end if;
  end process  Energy_Bin_950;    
  
  Energy_Bin_951 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_951   <=  (others =>'0');
		Energy_Bin_Rdy_951 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E951_C1_L and PEAK_C1 <= s_E951_C1_H and Bin_OR = '0') then
         s_Energy_Bin_951 <= s_Energy_Bin_951 +'1';
		 Energy_Bin_Rdy_951 <= '1';
		else
		 s_Energy_Bin_951 <= s_Energy_Bin_951;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_951 <= '0';
      end if;
    end if;
  end process  Energy_Bin_951;   
  
  Energy_Bin_952 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_952   <=  (others =>'0');
	    Energy_Bin_Rdy_952 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E952_C1_L and PEAK_C1 <= s_E952_C1_H and Bin_OR = '0') then
         s_Energy_Bin_952 <= s_Energy_Bin_952 +'1';
		 Energy_Bin_Rdy_952 <= '1';
		else
		 s_Energy_Bin_952 <= s_Energy_Bin_952;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_952 <= '0';
      end if;
    end if;
  end process  Energy_Bin_952;   
  
  Energy_Bin_953 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_953   <=  (others =>'0');
	    Energy_Bin_Rdy_953 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E953_C1_L and PEAK_C1 <= s_E953_C1_H and Bin_OR = '0') then
         s_Energy_Bin_953 <= s_Energy_Bin_953 +'1';
		 Energy_Bin_Rdy_953 <= '1';
		else
		 s_Energy_Bin_953 <= s_Energy_Bin_953;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_953 <= '0';
      end if;
    end if;
  end process  Energy_Bin_953;   
  
  Energy_Bin_954 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_954   <=  (others =>'0');
		Energy_Bin_Rdy_954 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E954_C1_L and PEAK_C1 <= s_E954_C1_H and Bin_OR = '0') then
         s_Energy_Bin_954 <= s_Energy_Bin_954 +'1';
		 Energy_Bin_Rdy_954 <= '1';
		else
		 s_Energy_Bin_954 <= s_Energy_Bin_954;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_954 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_954;   
 
 
  Energy_Bin_955 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_955   <=  (others =>'0');
		Energy_Bin_Rdy_955 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E955_C1_L and PEAK_C1 <= s_E955_C1_H and Bin_OR = '0') then
         s_Energy_Bin_955 <= s_Energy_Bin_955 +'1';
		 Energy_Bin_Rdy_955 <= '1';
		else
		 s_Energy_Bin_955 <= s_Energy_Bin_955;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_955 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_955;  
 
  
  Energy_Bin_956 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_956   <=  (others =>'0');
		Energy_Bin_Rdy_956 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E956_C1_L and PEAK_C1 <= s_E956_C1_H and Bin_OR = '0') then
         s_Energy_Bin_956 <= s_Energy_Bin_956 +'1';
		 Energy_Bin_Rdy_956 <= '1';
		else
		 s_Energy_Bin_956 <= s_Energy_Bin_956;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_956 <= '0';
      end if;
    end if;
  end process  Energy_Bin_956;   
  
 Energy_Bin_957 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_957   <=  (others =>'0');
		Energy_Bin_Rdy_957 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E957_C1_L and PEAK_C1 <= s_E957_C1_H and Bin_OR = '0') then
         s_Energy_Bin_957 <= s_Energy_Bin_957 +'1';
		 Energy_Bin_Rdy_957 <= '1';
		else
		 s_Energy_Bin_957 <= s_Energy_Bin_957;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_957 <= '0';
      end if;
    end if;
  end process  Energy_Bin_957;   
  
  Energy_Bin_958 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_958   <=  (others =>'0');
		Energy_Bin_Rdy_958 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E958_C1_L and PEAK_C1 <= s_E958_C1_H and Bin_OR = '0') then
         s_Energy_Bin_958 <= s_Energy_Bin_958 +'1';
		 Energy_Bin_Rdy_958 <= '1';
		else
		 s_Energy_Bin_958 <= s_Energy_Bin_958;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_958 <= '0';
      end if;
    end if;
  end process  Energy_Bin_958;   
  
  Energy_Bin_959 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_959   <=  (others =>'0');
		Energy_Bin_Rdy_959 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E959_C1_L and PEAK_C1 <= s_E959_C1_H and Bin_OR = '0') then
         s_Energy_Bin_959 <= s_Energy_Bin_959 +'1';
		 Energy_Bin_Rdy_959 <= '1';
		else
		 s_Energy_Bin_959 <= s_Energy_Bin_959;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_959 <= '0';
      end if;
    end if;
  end process  Energy_Bin_959;           
  
     Energy_Bin_960 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_960   <=  (others =>'0');
		Energy_Bin_Rdy_960 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E960_C1_L and PEAK_C1 <= s_E960_C1_H and Bin_OR = '0') then
         s_Energy_Bin_960 <= s_Energy_Bin_960 +'1';
		 Energy_Bin_Rdy_960 <= '1';
		else
		 s_Energy_Bin_960 <= s_Energy_Bin_960;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_960 <= '0';
      end if;
    end if;
  end process  Energy_Bin_960;    
  
  Energy_Bin_961 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_961   <=  (others =>'0');
		Energy_Bin_Rdy_961 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E961_C1_L and PEAK_C1 <= s_E961_C1_H and Bin_OR = '0') then
         s_Energy_Bin_961 <= s_Energy_Bin_961 +'1';
		 Energy_Bin_Rdy_961 <= '1';
		else
		 s_Energy_Bin_961 <= s_Energy_Bin_961;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_961 <= '0';
      end if;
    end if;
  end process  Energy_Bin_961;   
  
  Energy_Bin_962 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_962   <=  (others =>'0');
	    Energy_Bin_Rdy_962 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E962_C1_L and PEAK_C1 <= s_E962_C1_H and Bin_OR = '0') then
         s_Energy_Bin_962 <= s_Energy_Bin_962 +'1';
		 Energy_Bin_Rdy_962 <= '1';
		else
		 s_Energy_Bin_962 <= s_Energy_Bin_962;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_962 <= '0';
      end if;
    end if;
  end process  Energy_Bin_962;   
  
  Energy_Bin_963 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_963   <=  (others =>'0');
	    Energy_Bin_Rdy_963 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E963_C1_L and PEAK_C1 <= s_E963_C1_H and Bin_OR = '0') then
         s_Energy_Bin_963 <= s_Energy_Bin_963 +'1';
		 Energy_Bin_Rdy_963 <= '1';
		else
		 s_Energy_Bin_963 <= s_Energy_Bin_963;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_963 <= '0';
      end if;
    end if;
  end process  Energy_Bin_963;   
  
  Energy_Bin_964 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_964   <=  (others =>'0');
		Energy_Bin_Rdy_964 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E964_C1_L and PEAK_C1 <= s_E964_C1_H and Bin_OR = '0') then
         s_Energy_Bin_964 <= s_Energy_Bin_964 +'1';
		 Energy_Bin_Rdy_964 <= '1';
		else
		 s_Energy_Bin_964 <= s_Energy_Bin_964;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_964 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_964;   
 
 
  Energy_Bin_965 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_965   <=  (others =>'0');
		Energy_Bin_Rdy_965 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E965_C1_L and PEAK_C1 <= s_E965_C1_H and Bin_OR = '0') then
         s_Energy_Bin_965 <= s_Energy_Bin_965 +'1';
		 Energy_Bin_Rdy_965 <= '1';
		else
		 s_Energy_Bin_965 <= s_Energy_Bin_965;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_965 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_965;  
 
  
  Energy_Bin_966 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_966   <=  (others =>'0');
		Energy_Bin_Rdy_966 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E966_C1_L and PEAK_C1 <= s_E966_C1_H and Bin_OR = '0') then
         s_Energy_Bin_966 <= s_Energy_Bin_966 +'1';
		 Energy_Bin_Rdy_966 <= '1';
		else
		 s_Energy_Bin_966 <= s_Energy_Bin_966;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_966 <= '0';
      end if;
    end if;
  end process  Energy_Bin_966;   
  
 Energy_Bin_967 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_967   <=  (others =>'0');
		Energy_Bin_Rdy_967 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E967_C1_L and PEAK_C1 <= s_E967_C1_H and Bin_OR = '0') then
         s_Energy_Bin_967 <= s_Energy_Bin_967 +'1';
		 Energy_Bin_Rdy_967 <= '1';
		else
		 s_Energy_Bin_967 <= s_Energy_Bin_967;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_967 <= '0';
      end if;
    end if;
  end process  Energy_Bin_967;   
  
  Energy_Bin_968 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_968   <=  (others =>'0');
		Energy_Bin_Rdy_968 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E968_C1_L and PEAK_C1 <= s_E968_C1_H and Bin_OR = '0') then
         s_Energy_Bin_968 <= s_Energy_Bin_968 +'1';
		 Energy_Bin_Rdy_968 <= '1';
		else
		 s_Energy_Bin_968 <= s_Energy_Bin_968;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_968 <= '0';
      end if;
    end if;
  end process  Energy_Bin_968;   
  
  Energy_Bin_969 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_969   <=  (others =>'0');
		Energy_Bin_Rdy_969 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E969_C1_L and PEAK_C1 <= s_E969_C1_H and Bin_OR = '0') then
         s_Energy_Bin_969 <= s_Energy_Bin_969 +'1';
		 Energy_Bin_Rdy_969 <= '1';
		else
		 s_Energy_Bin_969 <= s_Energy_Bin_969;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_969 <= '0';
      end if;
    end if;
  end process  Energy_Bin_969;         
  
     Energy_Bin_970 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_970   <=  (others =>'0');
		Energy_Bin_Rdy_970 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E970_C1_L and PEAK_C1 <= s_E970_C1_H and Bin_OR = '0') then
         s_Energy_Bin_970 <= s_Energy_Bin_970 +'1';
		 Energy_Bin_Rdy_970 <= '1';
		else
		 s_Energy_Bin_970 <= s_Energy_Bin_970;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_970 <= '0';
      end if;
    end if;
  end process  Energy_Bin_970;    
  
  Energy_Bin_971 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_971   <=  (others =>'0');
		Energy_Bin_Rdy_971 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E971_C1_L and PEAK_C1 <= s_E971_C1_H and Bin_OR = '0') then
         s_Energy_Bin_971 <= s_Energy_Bin_971 +'1';
		 Energy_Bin_Rdy_971 <= '1';
		else
		 s_Energy_Bin_971 <= s_Energy_Bin_971;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_971 <= '0';
      end if;
    end if;
  end process  Energy_Bin_971;   
  
  Energy_Bin_972 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_972   <=  (others =>'0');
	    Energy_Bin_Rdy_972 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E972_C1_L and PEAK_C1 <= s_E972_C1_H and Bin_OR = '0') then
         s_Energy_Bin_972 <= s_Energy_Bin_972 +'1';
		 Energy_Bin_Rdy_972 <= '1';
		else
		 s_Energy_Bin_972 <= s_Energy_Bin_972;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_972 <= '0';
      end if;
    end if;
  end process  Energy_Bin_972;   
  
  Energy_Bin_973 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_973   <=  (others =>'0');
	    Energy_Bin_Rdy_973 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E973_C1_L and PEAK_C1 <= s_E973_C1_H and Bin_OR = '0') then
         s_Energy_Bin_973 <= s_Energy_Bin_973 +'1';
		 Energy_Bin_Rdy_973 <= '1';
		else
		 s_Energy_Bin_973 <= s_Energy_Bin_973;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_973 <= '0';
      end if;
    end if;
  end process  Energy_Bin_973;   
  
  Energy_Bin_974 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_974   <=  (others =>'0');
		Energy_Bin_Rdy_974 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E974_C1_L and PEAK_C1 <= s_E974_C1_H and Bin_OR = '0') then
         s_Energy_Bin_974 <= s_Energy_Bin_974 +'1';
		 Energy_Bin_Rdy_974 <= '1';
		else
		 s_Energy_Bin_974 <= s_Energy_Bin_974;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_974 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_974;   
 
 
  Energy_Bin_975 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_975   <=  (others =>'0');
		Energy_Bin_Rdy_975 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E975_C1_L and PEAK_C1 <= s_E975_C1_H and Bin_OR = '0') then
         s_Energy_Bin_975 <= s_Energy_Bin_975 +'1';
		 Energy_Bin_Rdy_975 <= '1';
		else
		 s_Energy_Bin_975 <= s_Energy_Bin_975;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_975 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_975;  
 
  
  Energy_Bin_976 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_976   <=  (others =>'0');
		Energy_Bin_Rdy_976 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E976_C1_L and PEAK_C1 <= s_E976_C1_H and Bin_OR = '0') then
         s_Energy_Bin_976 <= s_Energy_Bin_976 +'1';
		 Energy_Bin_Rdy_976 <= '1';
		else
		 s_Energy_Bin_976 <= s_Energy_Bin_976;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_976 <= '0';
      end if;
    end if;
  end process  Energy_Bin_976;   
  
 Energy_Bin_977 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_977   <=  (others =>'0');
		Energy_Bin_Rdy_977 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E977_C1_L and PEAK_C1 <= s_E977_C1_H and Bin_OR = '0') then
         s_Energy_Bin_977 <= s_Energy_Bin_977 +'1';
		 Energy_Bin_Rdy_977 <= '1';
		else
		 s_Energy_Bin_977 <= s_Energy_Bin_977;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_977 <= '0';
      end if;
    end if;
  end process  Energy_Bin_977;   
  
  Energy_Bin_978 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_978   <=  (others =>'0');
		Energy_Bin_Rdy_978 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E978_C1_L and PEAK_C1 <= s_E978_C1_H and Bin_OR = '0') then
         s_Energy_Bin_978 <= s_Energy_Bin_978 +'1';
		 Energy_Bin_Rdy_978 <= '1';
		else
		 s_Energy_Bin_978 <= s_Energy_Bin_978;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_978 <= '0';
      end if;
    end if;
  end process  Energy_Bin_978;   
  
  Energy_Bin_979 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_979   <=  (others =>'0');
		Energy_Bin_Rdy_979 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E979_C1_L and PEAK_C1 <= s_E979_C1_H and Bin_OR = '0') then
         s_Energy_Bin_979 <= s_Energy_Bin_979 +'1';
		 Energy_Bin_Rdy_979 <= '1';
		else
		 s_Energy_Bin_979 <= s_Energy_Bin_979;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_979 <= '0';
      end if;
    end if;
  end process  Energy_Bin_979;       
  
     Energy_Bin_980 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_980   <=  (others =>'0');
		Energy_Bin_Rdy_980 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E980_C1_L and PEAK_C1 <= s_E980_C1_H and Bin_OR = '0') then
         s_Energy_Bin_980 <= s_Energy_Bin_980 +'1';
		 Energy_Bin_Rdy_980 <= '1';
		else
		 s_Energy_Bin_980 <= s_Energy_Bin_980;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_980 <= '0';
      end if;
    end if;
  end process  Energy_Bin_980;    
  
  Energy_Bin_981 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_981   <=  (others =>'0');
		Energy_Bin_Rdy_981 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E981_C1_L and PEAK_C1 <= s_E981_C1_H and Bin_OR = '0') then
         s_Energy_Bin_981 <= s_Energy_Bin_981 +'1';
		 Energy_Bin_Rdy_981 <= '1';
		else
		 s_Energy_Bin_981 <= s_Energy_Bin_981;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_981 <= '0';
      end if;
    end if;
  end process  Energy_Bin_981;   
  
  Energy_Bin_982 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_982   <=  (others =>'0');
	    Energy_Bin_Rdy_982 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E982_C1_L and PEAK_C1 <= s_E982_C1_H and Bin_OR = '0') then
         s_Energy_Bin_982 <= s_Energy_Bin_982 +'1';
		 Energy_Bin_Rdy_982 <= '1';
		else
		 s_Energy_Bin_982 <= s_Energy_Bin_982;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_982 <= '0';
      end if;
    end if;
  end process  Energy_Bin_982;   
  
  Energy_Bin_983 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_983   <=  (others =>'0');
	    Energy_Bin_Rdy_983 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E983_C1_L and PEAK_C1 <= s_E983_C1_H and Bin_OR = '0') then
         s_Energy_Bin_983 <= s_Energy_Bin_983 +'1';
		 Energy_Bin_Rdy_983 <= '1';
		else
		 s_Energy_Bin_983 <= s_Energy_Bin_983;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_983 <= '0';
      end if;
    end if;
  end process  Energy_Bin_983;   
  
  Energy_Bin_984 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_984   <=  (others =>'0');
		Energy_Bin_Rdy_984 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E984_C1_L and PEAK_C1 <= s_E984_C1_H and Bin_OR = '0') then
         s_Energy_Bin_984 <= s_Energy_Bin_984 +'1';
		 Energy_Bin_Rdy_984 <= '1';
		else
		 s_Energy_Bin_984 <= s_Energy_Bin_984;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_984 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_984;   
 
 
  Energy_Bin_985 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_985   <=  (others =>'0');
		Energy_Bin_Rdy_985 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E985_C1_L and PEAK_C1 <= s_E985_C1_H and Bin_OR = '0') then
         s_Energy_Bin_985 <= s_Energy_Bin_985 +'1';
		 Energy_Bin_Rdy_985 <= '1';
		else
		 s_Energy_Bin_985 <= s_Energy_Bin_985;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_985 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_985;  
 
  
  Energy_Bin_986 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_986   <=  (others =>'0');
		Energy_Bin_Rdy_986 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E986_C1_L and PEAK_C1 <= s_E986_C1_H and Bin_OR = '0') then
         s_Energy_Bin_986 <= s_Energy_Bin_986 +'1';
		 Energy_Bin_Rdy_986 <= '1';
		else
		 s_Energy_Bin_986 <= s_Energy_Bin_986;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_986 <= '0';
      end if;
    end if;
  end process  Energy_Bin_986;   
  
 Energy_Bin_987 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_987   <=  (others =>'0');
		Energy_Bin_Rdy_987 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E987_C1_L and PEAK_C1 <= s_E987_C1_H and Bin_OR = '0') then
         s_Energy_Bin_987 <= s_Energy_Bin_987 +'1';
		 Energy_Bin_Rdy_987 <= '1';
		else
		 s_Energy_Bin_987 <= s_Energy_Bin_987;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_987 <= '0';
      end if;
    end if;
  end process  Energy_Bin_987;   
  
  Energy_Bin_988 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_988   <=  (others =>'0');
		Energy_Bin_Rdy_988 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E988_C1_L and PEAK_C1 <= s_E988_C1_H and Bin_OR = '0') then
         s_Energy_Bin_988 <= s_Energy_Bin_988 +'1';
		 Energy_Bin_Rdy_988 <= '1';
		else
		 s_Energy_Bin_988 <= s_Energy_Bin_988;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_988 <= '0';
      end if;
    end if;
  end process  Energy_Bin_988;   
  
  Energy_Bin_989 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_989   <=  (others =>'0');
		Energy_Bin_Rdy_989 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E989_C1_L and PEAK_C1 <= s_E989_C1_H and Bin_OR = '0') then
         s_Energy_Bin_989 <= s_Energy_Bin_989 +'1';
		 Energy_Bin_Rdy_989 <= '1';
		else
		 s_Energy_Bin_989 <= s_Energy_Bin_989;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_989 <= '0';
      end if;
    end if;
  end process  Energy_Bin_989;      
  
     Energy_Bin_990 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_990   <=  (others =>'0');
		Energy_Bin_Rdy_990 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E990_C1_L and PEAK_C1 <= s_E990_C1_H and Bin_OR = '0') then
         s_Energy_Bin_990 <= s_Energy_Bin_990 +'1';
		 Energy_Bin_Rdy_990 <= '1';
		else
		 s_Energy_Bin_990 <= s_Energy_Bin_990;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_990 <= '0';
      end if;
    end if;
  end process  Energy_Bin_990;    
  
  Energy_Bin_991 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_991   <=  (others =>'0');
		Energy_Bin_Rdy_991 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E991_C1_L and PEAK_C1 <= s_E991_C1_H and Bin_OR = '0') then
         s_Energy_Bin_991 <= s_Energy_Bin_991 +'1';
		 Energy_Bin_Rdy_991 <= '1';
		else
		 s_Energy_Bin_991 <= s_Energy_Bin_991;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_991 <= '0';
      end if;
    end if;
  end process  Energy_Bin_991;   
  
  Energy_Bin_992 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_992   <=  (others =>'0');
	    Energy_Bin_Rdy_992 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E992_C1_L and PEAK_C1 <= s_E992_C1_H and Bin_OR = '0') then
         s_Energy_Bin_992 <= s_Energy_Bin_992 +'1';
		 Energy_Bin_Rdy_992 <= '1';
		else
		 s_Energy_Bin_992 <= s_Energy_Bin_992;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_992 <= '0';
      end if;
    end if;
  end process  Energy_Bin_992;   
  
  Energy_Bin_993 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_993   <=  (others =>'0');
	    Energy_Bin_Rdy_993 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E993_C1_L and PEAK_C1 <= s_E993_C1_H and Bin_OR = '0') then
         s_Energy_Bin_993 <= s_Energy_Bin_993 +'1';
		 Energy_Bin_Rdy_993 <= '1';
		else
		 s_Energy_Bin_993 <= s_Energy_Bin_993;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_993 <= '0';
      end if;
    end if;
  end process  Energy_Bin_993;   
  
  Energy_Bin_994 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_994   <=  (others =>'0');
		Energy_Bin_Rdy_994 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E994_C1_L and PEAK_C1 <= s_E994_C1_H and Bin_OR = '0') then
         s_Energy_Bin_994 <= s_Energy_Bin_994 +'1';
		 Energy_Bin_Rdy_994 <= '1';
		else
		 s_Energy_Bin_994 <= s_Energy_Bin_994;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_994 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_994;   
 
 
  Energy_Bin_995 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_995   <=  (others =>'0');
		Energy_Bin_Rdy_995 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E995_C1_L and PEAK_C1 <= s_E995_C1_H and Bin_OR = '0') then
         s_Energy_Bin_995 <= s_Energy_Bin_995 +'1';
		 Energy_Bin_Rdy_995 <= '1';
		else
		 s_Energy_Bin_995 <= s_Energy_Bin_995;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_995 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_995;  
 
  
  Energy_Bin_996 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_996   <=  (others =>'0');
		Energy_Bin_Rdy_996 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E996_C1_L and PEAK_C1 <= s_E996_C1_H and Bin_OR = '0') then
         s_Energy_Bin_996 <= s_Energy_Bin_996 +'1';
		 Energy_Bin_Rdy_996 <= '1';
		else
		 s_Energy_Bin_996 <= s_Energy_Bin_996;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_996 <= '0';
      end if;
    end if;
  end process  Energy_Bin_996;   
  
 Energy_Bin_997 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_997   <=  (others =>'0');
		Energy_Bin_Rdy_997 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E997_C1_L and PEAK_C1 <= s_E997_C1_H and Bin_OR = '0') then
         s_Energy_Bin_997 <= s_Energy_Bin_997 +'1';
		 Energy_Bin_Rdy_997 <= '1';
		else
		 s_Energy_Bin_997 <= s_Energy_Bin_997;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_997 <= '0';
      end if;
    end if;
  end process  Energy_Bin_997;   
  
  Energy_Bin_998 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_998   <=  (others =>'0');
		Energy_Bin_Rdy_998 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E998_C1_L and PEAK_C1 <= s_E998_C1_H and Bin_OR = '0') then
         s_Energy_Bin_998 <= s_Energy_Bin_998 +'1';
		 Energy_Bin_Rdy_998 <= '1';
		else
		 s_Energy_Bin_998 <= s_Energy_Bin_998;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_998 <= '0';
      end if;
    end if;
  end process  Energy_Bin_998;   
  
  Energy_Bin_999 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_999   <=  (others =>'0');
		Energy_Bin_Rdy_999 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E999_C1_L and PEAK_C1 <= s_E999_C1_H and Bin_OR = '0') then
         s_Energy_Bin_999 <= s_Energy_Bin_999 +'1';
		 Energy_Bin_Rdy_999 <= '1';
		else
		 s_Energy_Bin_999 <= s_Energy_Bin_999;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_999 <= '0';
      end if;
    end if;
  end process  Energy_Bin_999;   

    Energy_Bin_1000 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1000   <=  (others =>'0');
		Energy_Bin_Rdy_1000 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E1000_C1_L and PEAK_C1 <= s_E1000_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1000 <= s_Energy_Bin_1000 +'1';
		 Energy_Bin_Rdy_1000 <= '1';
		else
		 s_Energy_Bin_1000 <= s_Energy_Bin_1000;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1000 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1000;    
  
  Energy_Bin_1001 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1001   <=  (others =>'0');
		Energy_Bin_Rdy_1001 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E1001_C1_L and PEAK_C1 <= s_E1001_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1001 <= s_Energy_Bin_1001 +'1';
		 Energy_Bin_Rdy_1001 <= '1';
		else
		 s_Energy_Bin_1001 <= s_Energy_Bin_1001;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1001 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1001;   
  
  Energy_Bin_1002 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1002   <=  (others =>'0');
	    Energy_Bin_Rdy_1002 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E1002_C1_L and PEAK_C1 <= s_E1002_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1002 <= s_Energy_Bin_1002 +'1';
		 Energy_Bin_Rdy_1002 <= '1';
		else
		 s_Energy_Bin_1002 <= s_Energy_Bin_1002;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1002 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1002;   
  
  Energy_Bin_1003 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1003   <=  (others =>'0');
	    Energy_Bin_Rdy_1003 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E1003_C1_L and PEAK_C1 <= s_E1003_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1003 <= s_Energy_Bin_1003 +'1';
		 Energy_Bin_Rdy_1003 <= '1';
		else
		 s_Energy_Bin_1003 <= s_Energy_Bin_1003;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1003 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1003;   
  
  Energy_Bin_1004 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1004   <=  (others =>'0');
		Energy_Bin_Rdy_1004 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E1004_C1_L and PEAK_C1 <= s_E1004_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1004 <= s_Energy_Bin_1004 +'1';
		 Energy_Bin_Rdy_1004 <= '1';
		else
		 s_Energy_Bin_1004 <= s_Energy_Bin_1004;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1004 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_1004;   
 
 
  Energy_Bin_1005 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1005   <=  (others =>'0');
		Energy_Bin_Rdy_1005 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E1005_C1_L and PEAK_C1 <= s_E1005_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1005 <= s_Energy_Bin_1005 +'1';
		 Energy_Bin_Rdy_1005 <= '1';
		else
		 s_Energy_Bin_1005 <= s_Energy_Bin_1005;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1005 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_1005;  
 
  
  Energy_Bin_1006 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1006   <=  (others =>'0');
		Energy_Bin_Rdy_1006 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E1006_C1_L and PEAK_C1 <= s_E1006_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1006 <= s_Energy_Bin_1006 +'1';
		 Energy_Bin_Rdy_1006 <= '1';
		else
		 s_Energy_Bin_1006 <= s_Energy_Bin_1006;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1006 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1006;   
  
 Energy_Bin_1007 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1007   <=  (others =>'0');
		Energy_Bin_Rdy_1007 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E1007_C1_L and PEAK_C1 <= s_E1007_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1007 <= s_Energy_Bin_1007 +'1';
		 Energy_Bin_Rdy_1007 <= '1';
		else
		 s_Energy_Bin_1007 <= s_Energy_Bin_1007;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1007 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1007;   
  
  Energy_Bin_1008 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1008   <=  (others =>'0');
		Energy_Bin_Rdy_1008 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E1008_C1_L and PEAK_C1 <= s_E1008_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1008 <= s_Energy_Bin_1008 +'1';
		 Energy_Bin_Rdy_1008 <= '1';
		else
		 s_Energy_Bin_1008 <= s_Energy_Bin_1008;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1008 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1008;   
  
  Energy_Bin_1009 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1009   <=  (others =>'0');
		Energy_Bin_Rdy_1009 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E1009_C1_L and PEAK_C1 <= s_E1009_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1009 <= s_Energy_Bin_1009 +'1';
		 Energy_Bin_Rdy_1009 <= '1';
		else
		 s_Energy_Bin_1009 <= s_Energy_Bin_1009;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1009 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1009;      
  
     Energy_Bin_1010 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1010   <=  (others =>'0');
		Energy_Bin_Rdy_1010 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E1010_C1_L and PEAK_C1 <= s_E1010_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1010 <= s_Energy_Bin_1010 +'1';
		 Energy_Bin_Rdy_1010 <= '1';
		else
		 s_Energy_Bin_1010 <= s_Energy_Bin_1010;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1010 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1010;    
  
  Energy_Bin_1011 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1011   <=  (others =>'0');
		Energy_Bin_Rdy_1011 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E1011_C1_L and PEAK_C1 <= s_E1011_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1011 <= s_Energy_Bin_1011 +'1';
		 Energy_Bin_Rdy_1011 <= '1';
		else
		 s_Energy_Bin_1011 <= s_Energy_Bin_1011;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1011 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1011;   
  
  Energy_Bin_1012 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1012   <=  (others =>'0');
	    Energy_Bin_Rdy_1012 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E1012_C1_L and PEAK_C1 <= s_E1012_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1012 <= s_Energy_Bin_1012 +'1';
		 Energy_Bin_Rdy_1012 <= '1';
		else
		 s_Energy_Bin_1012 <= s_Energy_Bin_1012;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1012 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1012;   
  
  Energy_Bin_1013 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1013   <=  (others =>'0');
	    Energy_Bin_Rdy_1013 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E1013_C1_L and PEAK_C1 <= s_E1013_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1013 <= s_Energy_Bin_1013 +'1';
		 Energy_Bin_Rdy_1013 <= '1';
		else
		 s_Energy_Bin_1013 <= s_Energy_Bin_1013;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1013 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1013;   
  
  Energy_Bin_1014 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1014   <=  (others =>'0');
		Energy_Bin_Rdy_1014 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E1014_C1_L and PEAK_C1 <= s_E1014_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1014 <= s_Energy_Bin_1014 +'1';
		 Energy_Bin_Rdy_1014 <= '1';
		else
		 s_Energy_Bin_1014 <= s_Energy_Bin_1014;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1014 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_1014;   
 
 
  Energy_Bin_1015 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1015   <=  (others =>'0');
		Energy_Bin_Rdy_1015 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E1015_C1_L and PEAK_C1 <= s_E1015_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1015 <= s_Energy_Bin_1015 +'1';
		 Energy_Bin_Rdy_1015 <= '1';
		else
		 s_Energy_Bin_1015 <= s_Energy_Bin_1015;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1015 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_1015;  
 
  
  Energy_Bin_1016 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1016   <=  (others =>'0');
		Energy_Bin_Rdy_1016 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E1016_C1_L and PEAK_C1 <= s_E1016_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1016 <= s_Energy_Bin_1016 +'1';
		 Energy_Bin_Rdy_1016 <= '1';
		else
		 s_Energy_Bin_1016 <= s_Energy_Bin_1016;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1016 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1016;   
  
 Energy_Bin_1017 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1017   <=  (others =>'0');
		Energy_Bin_Rdy_1017 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E1017_C1_L and PEAK_C1 <= s_E1017_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1017 <= s_Energy_Bin_1017 +'1';
		 Energy_Bin_Rdy_1017 <= '1';
		else
		 s_Energy_Bin_1017 <= s_Energy_Bin_1017;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1017 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1017;   
  
  Energy_Bin_1018 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1018   <=  (others =>'0');
		Energy_Bin_Rdy_1018 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E1018_C1_L and PEAK_C1 <= s_E1018_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1018 <= s_Energy_Bin_1018 +'1';
		 Energy_Bin_Rdy_1018 <= '1';
		else
		 s_Energy_Bin_1018 <= s_Energy_Bin_1018;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1018 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1018;   
  
  Energy_Bin_1019 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1019   <=  (others =>'0');
		Energy_Bin_Rdy_1019 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E1019_C1_L and PEAK_C1 <= s_E1019_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1019 <= s_Energy_Bin_1019 +'1';
		 Energy_Bin_Rdy_1019 <= '1';
		else
		 s_Energy_Bin_1019 <= s_Energy_Bin_1019;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1019 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1019;       
  
     Energy_Bin_1020 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1020   <=  (others =>'0');
		Energy_Bin_Rdy_1020 <= '0';
      elsif(PEAK_FL_Ris = '1' ) then
	  
	    if(PEAK_C1 > s_E1020_C1_L and PEAK_C1 <= s_E1020_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1020 <= s_Energy_Bin_1020 +'1';
		 Energy_Bin_Rdy_1020 <= '1';
		else
		 s_Energy_Bin_1020 <= s_Energy_Bin_1020;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1020 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1020;    
  
  Energy_Bin_1021 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1021   <=  (others =>'0');
		Energy_Bin_Rdy_1021 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E1021_C1_L and PEAK_C1 <= s_E1021_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1021 <= s_Energy_Bin_1021 +'1';
		 Energy_Bin_Rdy_1021 <= '1';
		else
		 s_Energy_Bin_1021 <= s_Energy_Bin_1021;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1021 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1021;   
  
  Energy_Bin_1022 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1022   <=  (others =>'0');
	    Energy_Bin_Rdy_1022 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E1022_C1_L and PEAK_C1 <= s_E1022_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1022 <= s_Energy_Bin_1022 +'1';
		 Energy_Bin_Rdy_1022 <= '1';
		else
		 s_Energy_Bin_1022 <= s_Energy_Bin_1022;
		end if;
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1022 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1022;   
  
  Energy_Bin_1023 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1023   <=  (others =>'0');
	    Energy_Bin_Rdy_1023 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E1023_C1_L and PEAK_C1 <= s_E1023_C1_H and Bin_OR = '0') then
         s_Energy_Bin_1023 <= s_Energy_Bin_1023 +'1';
		 Energy_Bin_Rdy_1023 <= '1';
		else
		 s_Energy_Bin_1023 <= s_Energy_Bin_1023;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1023 <= '0';
      end if;
    end if;
  end process  Energy_Bin_1023;   
  
  Energy_Bin_1024 : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_1024   <=  (others =>'0');
		Energy_Bin_Rdy_1024 <= '0';
      elsif(PEAK_FL_Ris = '1') then
	  
	    if(PEAK_C1 > s_E1024_C1_L and PEAK_C1 < s_E1024_C1_H and Bin_OR = '0') then -- ************************************************************************** S_E1024_c1_H = 2048; PEAK_C1 < s_E1024_C1_H.
         s_Energy_Bin_1024 <= s_Energy_Bin_1024 +'1';
		 Energy_Bin_Rdy_1024 <= '1';
		else
		 s_Energy_Bin_1024 <= s_Energy_Bin_1024;
		end if;
		
	  elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_1024 <= '0';
      
      end if;
    end if;
  end process  Energy_Bin_1024;   


  Energy_Bin_reject : process (CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        s_Energy_Bin_reject   <=  (others =>'0');
        Energy_Bin_Rdy_reject <= '0';
      elsif(PEAK_FL_Ris_s = '1' ) then
	    if(Energy_Bin_Rdy = '0') then
         s_Energy_Bin_reject <= s_Energy_Bin_reject +'1';
         Energy_Bin_Rdy_reject <= '1';
		else
		 s_Energy_Bin_reject <= s_Energy_Bin_reject;
		end if;
		
      elsif(Energy_Ris_Dis = '1') then
	    Energy_Bin_Rdy_reject <= '0';
      end if;
    end if;
 end process  Energy_Bin_reject;    
  
/*   Energy_Bin_REG_OR_det : process(CLK100)
  begin
    if (rising_edge(CLK100))then
      if (RST = '1') then
        Bin_OR <= '0';  
      elsif(s_Energy_Bin_1 < x"FFFFFFFD" and s_Energy_Bin_2 < x"FFFFFFFD" and s_Energy_Bin_3 < x"FFFFFFFD" and s_Energy_Bin_4 < x"FFFFFFFD" and s_Energy_Bin_5 < x"FFFFFFFD" and s_Energy_Bin_6 < x"FFFFFFFD" and s_Energy_Bin_7 < x"FFFFFFFD" and s_Energy_Bin_8 < x"FFFFFFFD" and s_Energy_Bin_9 < x"FFFFFFFD" and s_Energy_Bin_10 < x"FFFFFFFD") then 
        Bin_OR <= '0';
      else
        Bin_OR <= '1';
      end if;
    end if;
  end process  Energy_Bin_REG_OR_det;   */
  
end architecture PeakDetector_RTL;
--============================================================================
-- Architecture definition section end - RTL
--****************************************************************************


--****************************************************************************
-- Module trailer section starts
--============================================================================
--
--
--
--
--
--============================================================================
-- Module trailer section ends
--****************************************************************************